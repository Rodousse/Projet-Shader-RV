MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���3�`�`�`��`锃`�� `���`�R�`�`�`���`��`˔�`��`�`��`�`Rich�`                PE  L �0N        � !	  �  �      �3                               �                              �+ Y   �% (                            p `  `                            � @                                         .text   %�     �                   `.rdata  I,      .   �             @  @.data   1   0                   @  �.reloc  �$   p  &   6             @  B                                                                                                                                                                                                                                                                                                                                                                                                        U��E��dt���   uB��D    ]á�D�H�Q8��+�D=�  |�&  ��D�H�Q8�ң�D�   ]��������U�졨D�UV��H�ApVR�Ѓ���^]� ��������������U�졨DV��H�Q`V�ҡ�D�H�U�ApVR�Ѓ���^]� U�졨DV��H�Q`V�ҡ�D�U�H�E�IdRj�PV�у���^]� ����������U�졨DVW�}��H�Q`W�ҡ�D�H�U�E�I4RPV�ы�����t"��D�B�HpWV�ы�D�B�HV�у���_^]� ���������������U�졨DVW�}��H�Q`W�ҡ�D�H�QLV�ҋ�����t ��D�H�QpWV�ҡ�D�H�QV�҃���_^]� ���������U���,�EV�]�W�E3��]�3��E�]��3��U���  �E�E�M�E�P�M�Q�M��E�   �U��E�   �8  �U�R����;  ����u�E�PS�`A  ������t~V���<  ��D���   ���   jj���Ћ���tV��D���   �E�Rlj P���҅�t9��D�D�ԋ��   Q�$�ȋB0V�ЍM��~)  G���4���_�   ^��]ÍM��a)  _3�^��]����������U��QV�u���AJ  �E���t}���$    ���D���   �ȋB��=/  t)-�  t"���=��t��D���   �M��B(���'��D���   �M��BL�ЍM�Q�C  ������I  �E���u�^��]���������U��V�u��tB��I V�J�����D���   �B4������P�������D���   �B(�����Ћ���u�^]�U�졨D�H�A`�� S�U�VR�Ћ�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҍE�P�M�Q荂  ��D���B�Pl�M�Q���ҋu��$V��t@��D�H�Q`�ҡ�D�H�Qdj j�h�V�ҡ�D�H�Al�U�R�Ѓ���^[��]Ë�D�Q�B`�Ћ�D�Q�Jp�E�VP�ы�D�B�Pl�M�Q�҃���^[��]��������������U���0  �13ŉE�V�u����  ������Ph  �  ��t������Q���������  �������jR芖  ��P���_�  �������d�  �M���3�^�) ��]����U��Q����G  �E�����   ���$    ���D���   �ȋB�Ћ�D=L  uN�Q@�E��JhP�у�h�  ��蕰  ��u)��D���   �M��PL�ҍE�P�4A  �����ZG  ���D���   �M��B(�ЉE����y�����]������U��V�u��t>��I �;�����D���   �B4����P�������D���   �B(�����Ћ���u�3�^]����;�  P����Y����U���HSV�uW����  �}�]��    ����  ��D���   �Bx���Ћ�D���   �E�Bx���Ћ�D�Q�M�R j QP�҃����v  ��D���   �B����=  ��   ��D���   �B����=  ��   ��D�QH�J(�E�VP�ы�H�U�P��D�M��HH�A8�U��U�VR�Ћ�P�@�M��D�U�QH�J0�E��E�VP�ы�H�U܋P���ĉM��M��M��U�U�h�  �PW�H�9����U�M���ĉ�U�h�  �HW�P�����M܋U����ĉ�M�h�  �PW�H���������D���   �P4���ҋM�UWQRP��D���   �B4����P�O�����D���   �B(�����Ћ�D���   ���B(���Ћ؅��:���_^[��]����U�����D���   �SVW�}j j �������]������]���  P������]��;]�]r�E���]��{�  �E�E�M�Q���}����]����]����  �U�R�����  jjj ����  �E�PVW��蠱  P��蘱  P�b���C��;]�]~���M��]�Q�����]���  _��^[��]�����U�졨D�H�A�U��DR�Ѓ���u��D�Q�Jl�EP�у�3���]Ë�D�B�P`�M�Q�ҡ�D�H�A`�U�R�Ћ�D�Q���   ��j �E�Pj=�M�҅�u>��D�H�Al�U�R�Ћ�D�Q�Jl�E�P�ы�D�B�Pl�MQ�҃�3���]ËM�V�E�PQj �U�R�M��������e�����D�Q�Rp�M�QP�ҡ�D�H�Al�U�R�Ћ�D�Q�Jl�E�P�ы�D�B�P�MQ�ҋM�+���HPAQ�E�P�M������D�Q�Rp�M�QP�ҡ�D�H�Al�U�R�Ћ�D�Q�E�RpP�M�Q�ҡ�D�H�A`�U�R�Ћ�D�Qj j�h��E̋JdP�ы�D�B�@ j �M�Q�U�R�Ћ�D�Q�Jl���ލE��PF�у�8��tB��D�B�Pl�M�Q�ҡ�D�H�Al�U�R�Ћ�D�Q�Jl�EP�у��   ^��]�j h��M��f�����D�B�@ j �M�Q�U�R�Ћ�D�Q�Jl���ލE��PF�у���tB��D�B�Pl�M�Q�ҡ�D�H�Al�U�R�Ћ�D�Q�Jl�EP�у��   ^��]�j h��M�������U�R�M���  ��D�H�Al�U�R�Ѓ���tB��D�Q�Jl�E�P�ы�D�B�Pl�M�Q�ҡ�D�H�Al�UR�Ѓ��   ^��]�j h��M��f����M�Q�M��Z  ��D���B�Pl�M�Q�҃���tB��D�H�Al�U�R�Ћ�D�Q�Jl�E�P�ы�D�B�Pl�MQ�҃��   ^��]�j h��M�������E�P�M���  ��D�Q�Jl���E�P�ы�D�B�Pl�M܃�Q�ҡ�D�H�Al�U�R�Ћ�D�Q�Jl�EP�у���t
�   ^��]�3�^��]���������������U���   SVW3�9=0t3�0��I �0jV�u���  ���E���uBG�<�0 ��0u׍M��|  �M$��|  ��D�H�Al�U@R�Ѓ�_^�'  [��]Ê�0�]���tEj P�n�  ����u1�M�|  �M$�|  ��D�Q�Jl�E@P�у�_^�'  [��]Ë�D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�Ѓ��M�Q�M��}  ��D���B�Pl�M�Q�E��҃��}� �Mt-�"|  �M$�|  ��D�H�Al�U@R�Ѓ�_^�'  [��]�j jQ�E�    �	�  ���E��M��u.��{  �M$��{  ��D�B�Pl�M@Q�҃�_^�'  [��]ÍE�P�5�  �M�P�l�  �M��{  �M$�<|  ���  �M$Q�M�{  �M$��|  j h��M������U�R�M$��|  ��D�H�Al�U�R�Ѓ��M$j Q��  ����t�U$j R��  ���M��	�  P�s����M���舳  ��D3�����3����  �����E�������  �ۍ�	�  O��ۉMȊM����  ��K���%�  H�E������%�  H�E������%�  H�M��E�3��j�  ��D�u����   �P�M�Q�M�j�ҋE�����   ��D�Q@P�Bh�Ћ�������   j j �M�Q����  jh�  ���I�  jh�  ���;�  j h�  ���-�  �U�jR��� �  �E�j P����  j W���	�  ��Q�$S���k�  ��Q�M��$Q���V�  ���U�Q�$R���A�  ���E�Q�$P���,�  �EP�MT;�}Q�M�PQ�7������E���l���j	R�sd  �E�jP�hd  ���M�Q�M��  Pj	�d  ���M��Fy  ��D�B�P�M@Q�҃���t"�E@P�M���x  �M�Qj�Fd  ���M��y  �ŰM�Rj �E$PQ訾  ������tj j V�M��  ��l���Rj	�d  �E�Pj��c  �M�Q落  ���M��x  ��l����x  �M���  �M�x  �M$�x  ��D�B�Pl�M@Q�҃������_%����^'  [��]�j h��M��w����M�Q�M$��y  ��D���B�Pl�M�Q�E��҃��}� ������M�x  �M$�x  ��D�H�Al�U@R�Ѓ�_^�'  [��]�������U����  �{  �E��E�P������ ���Q�������D�B�P�M�Q�҃���uE�� ����w  ��D�H�Al�U�R�ЍM�Q�\{  ��D�E�    �B�Pl�MQ�҃���]á�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�hdP�эU�R�E�P�M�Q�  �� P�M���v  P�� ���R�����P�/y  ���M��w  ��D�Q�Jl�E�P�ы�D�B�Pl�M�Q�ҡ�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�hTP�эU�R�E�P�M�Q��  ��(P�M��7v  P�� ���R������P�x  ���M��xv  ��D�Q�Jl�E�P�ы�D�B�Pl�M�Q�ҡ�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�ыE��='  ��  ��  ����  WPhH��,�������j h<���������j h4��<����������D�:�EP�M�Q�]  ��P������WR��  ��P��,���P������Q�f]  ��D��PR������P�o�  ��P�����Q��D���R�8]  P��<���P������Q�  ��P��$���R�  ��P������P�  ��P��d���Q�t  ��P��4���R�d  ��P��T���P�T  ��P��t���Q�D  ��P������R�4  ��P�M�������D�H�Al������R�Ћ�D�Q�Jl��t���P�ы�D�B�Pl��T���Q�ҡ�D�H�Al��4���R�Ћ�D�Q�Jl��d���P�ы�D�B�Pl������Q�ҡ�D�H�Al��$���R�Ћ�D�Q�Jl������P�ы�D�B�Pl��D���Q�ҡ�D�H�Al������R�Ћ�D�Q�Jl������P�ы�D�B������Q�Pl�ҡ�D�H�Al�U�R�Ћ�D�Q�Jl��<���P�ы�D�B�Pl�����Q�ҡ�D�H�Al��,���R�Ѓ�@_��  j h�M�������D�Q�Rp�E�P�M�Q�ҡ�D�H�Al�U�R�Ѓ��  �������0  �$�d* j h���\����C�����\���Q�M��������D�B�Pl��\���Q�҃��A  j h���L���������L���P�M�������D�Q�Jl��L���P�у��  j hp��l����������l���R�M��X�����D�H�Al��l���R�Ѓ���   j hH��|���������|���Q�M�������D�B�Pl��|���Q�҃��   j h�M��O����E�P�M��������D�Q�Jl�E�P�у��V��D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�Ћ�D�Q�Rp�E�P�M�Q�ҡ�D�H�Al�U�R�Ѓ� ��D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҡ�D�H�Ip�UR�E�P�ы�D�B�Pl�M�Q�ҡ�D�E�    �H��H  j j h   �ҋ�Dj �E��Q�JTh   P�E�P�ыM���<h1D4ChCD4Cjj j������R�u  ��D�H�AP�U�j R�ЋM���PQ�M��u  �M��u  j�����R������P��  j ������Q�  �U�R�|�  ��D�H�Al�U�R�Ѓ��������p  ������p  �� ����wp  ��D�Q�Jl�E�P�эU�R�,t  ��D�E�    �H�Al�UR�Ѓ���]Ðk' �' �' $( b( ��������U����   VW��s  h1D4ChCD4Cjj j�MQ�ȉE���s  ��D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�Ћ�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҡ�D�H�A`��x���R�Ћ�D�Q�Jdj j���x���h�P�ы�D�B�P`�M�Q�ҡ�D�H�Ad��@j j��U�h�R�Ћ�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҡ�D�E� �H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�ы�D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�ЋM���L3���s  ����  j j�M�Q�M���r  �E�<
�  <�  �M��s  f�U�H;���D�H�A`���u  ��8���R�Ћ�D�Q�JhV��8���jP�ы�D�B�P�M�Q�ҋ�D�Q��8���Q�J0P�E�P�ы�D�B�Pl��8���Q�ҋ�D�Q��$�E�P�B`����V�Ћ�D�Q�Jp�E�VP�у��K�������wp�$�42 j h���������������R�M��K�����D�H�Al�����R�Ѓ��/�M�Q�M��!�M���E�P��x�����M�Q�M���M��U�R������D�H�A`��X���R�Ћ�D�Q�Jdj j���X���h�P�ы�D�B�@p�M�Q��X���R�Ћ�D�Q�Jl��X���P����  ��(���R�Ћ�D�Q�JhV��(���jP�ы�D�B�P�M�Q�ҋ�D�Q��(���Q�J0P�E�P�ы�D�B�Pl��(���Q�҃�$�h  ��D�Q�E�P�B`����V�Ћ�D�Q�Jp�E�VP�у������������   �$�L2 ��D�B�P`��H���Q�ҡ�D�H�Adj j���H���h�R�Ћ�D�Q�Rp�E�P��H���Q�ҡ�D�H�Al��H���R�Ѓ� �h��D�Q�Rp�E�P�M�Q���M�U��6��D�B�@p��x���Q�U�R���-��D�Q�Rp�E�P�M�Q����U���D�H�IpR�E�P�у���D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�Ћ�D�Q�Rp�E�P�M�Q�ҡ�D�H�Al�U�R�Ѓ� �M�G�3p  ;��a����M��#o  �Mj Q��y  ��D�B�P`��h���Q�ҡ�D�H�Adj j���h���h�R�Ћ�D�Q�J�E�P�у� ��uV��D�B�P`�M�Q�ҡ�D�H�Adj j��U�htR�Ћ�D�Q�Rp�E�P�M�Q�ҡ�D�H�Al�U�R�Ѓ� ��D�Q�J�E�P�у���uV��D�B�P`�M�Q�ҡ�D�H�Adj j��U�htR�Ћ�D�Q�Rp�E�P�M�Q�ҡ�D�H�Al�U�R�Ѓ� ��D�Q�J<�E�j P�ы�D���B�P<�M�j Q�ҋ�D����h���QVP�B�H`����V�ы�D�B�Pp��x���VQ�҃��E���P�
i  ���U���R��h  ��������D�H�Q`��D��V�ҡ�D�H�Ap��h���VR�Ѓ�W�4�����D�Q�Jl��h���P�ы�D�B�Pl�M�Q�ҡ�D�H�Al�U�R�Ћ�D�Q�Jl�E�P�ы�D�B�Pl�M�Q�ҡ�D�H�Al��x���R�Ћ�D�Q�Jl�E�P�ы�D�B�Pl�M�Q�ҍE�P�Wl  ��8�M�E�    �uh  _^��]ÍI �, .- 7- <- H- Q- r. �. �. �. / &/ ������������U���   SV�P�  ������  ��    ��D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�эU�R�KQ  ��D�H�Al�U�R�Ћ�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҡ�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�у�D�U�R�E�P��t���Q�����  ���!h  P�U�R�E�P�  ��P�M�Q�  P�P  ��D�B�M��PlQ�ҡ�D�H�Al�U�R�Ћ�D�Q�Jl�E�P�ы�D�B�Pl�M�Q�҃� ��t�����f  ��D�H�Al�U�R�Ѓ���蠵  P�M�Q覾  P� P  ��D�B�Pl�M�Q�ҡ�D���   �B(�����Ћ����o�����D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҍE�P�O  ��D�Q�Jl�E�P�ы�D�B�P`�M�Q�ҡ�D�H�Adj j��U�hxR�ЍM�Q�rO  ��D�B�Pl�M�Q�ҡ�D���   ���   ��j��jS��  ��D����  ��D���   ���   ��3��Ѕ���  W��    ��D���   ���   V���Ћ�D�Q�J`���E�P�ы�D�B�Pdj j��M�h�Q�ҍE�P��N  ��D�Q�Jl�E�P�ы�D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�Ћ�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�҃�D�E�P�M�Q��t���R���m�  ���e  P�E�P�M�Q�  ��P�U�R��  P�N  ��D�H�Al�U�R�Ћ�D�Q�Jl�E�P�ы�D�B�Pl�M�Q�ҡ�D�H�Al�U�R�Ѓ� ��t����Qd  ��D�Q�Jl�E�P�у�����  P�U�R��  P�M  ��D�H�Al�U�R�Ћ�D���   ���   ����F��;��R���_^[��]������������U��E���   P������M�Q�������D�B�P�M�Q�҃���u"�M��c  ��D�H�Al�U�R�Ѓ�3���]Ë�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҍE�P�M�Q�U�R�  �� P��|�����b  P�E�P�M�Q�Oe  ����|����!c  ��D�B�Pl�M�Q�ҡ�D�H�Al�U�R�Ћ�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�҃��E�P�M��c  P�M�Q�U�R�  P�L  ��D�H�Al�U�R�Ћ�D�Q�Jl�E�P�ы�D�B�Pl�M�Q�ҍE�j P�q  ��$��tZ��D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�ЍM�Q�K  ��D�B�Pl�M�Q�ҍE���P��a  ��������M��b  �M���a  ��D�Q�Jl�E�P�у�3���]���U�졨D�P�Ej PQ�J �у����@]� �������������U�졨D�H�A`���U�VR�Ћ�D�Q�M�Rp�E�PQ�ҡ�D�H�A�U�R�Ћ�D�Q�MQ�J0P�E�P�ы�D�B�u�H`V�ы�D�B�Pp�M�VQ�ҡ�D�H�Al�U�R�Ѓ�,��^��]����������̡�D� �����  ;��@����������U�졨D�����������  v3���]Ë@�P`�M�Q�ҡ�D�H�Adj j��U�hR�ЍM�Q�J  ��D�B�Pl�M�Q�ҡ�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�эU�R��I  ��D�H�Al�U�R�Ѓ�8�   ��]�����������������������������U�졨D� ���=�  v3�]ËE�� t��t-Vu�u������   ]ù�D��  �����]�����U��E��D� ]�̡�D���   ���   �� Q��Y��������h�DPhD �0�  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h�DjhD �\�  ����t
�@��t]��3�]��������Vh�Dj\hD ���,�  ����t�@\��tV�Ѓ���^�����Vh�Dj`hD �����  ����t�@`��tV�Ѓ�^�������U��Vh�DjdhD �����  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�DjhhD ����  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�DjlhD ���L�  ����t�@l��tV�Ѓ�^�������U��Vh�Dh�   hD ����  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�Dh�   hD �����  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�DjphD ���y�  ����t�@p��t�MQV�Ѓ�^]� ��D^]� ��U��Vh�DjxhD ���9�  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�DjxhD �����  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�DjxhD ����  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������h�DjhD �_�  ����t	�@��t��3��������������U��V�u�> t+h�DjhD �#�  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h�DjhD ���  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�DjhD ����  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�DjhD ���Y�  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�Dj hD ����  ����t�@ ��tV�Ѓ�^�3�^���Vh�Dj$hD �����  ����t�@$��tV�Ѓ�^�3�^���U��Vh�Dj(hD ����  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�Dj,hD ���i�  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�Dj(hD ���)�  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�Dj4hD �����  ����t�@4��tV�Ѓ�^�3�^���U��Vh�Dj8hD ����  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�Dj<hD ���Y�  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�DjDhD ����  ����t�@D��tV�Ѓ�^�3�^���U��Vh�DjHhD �����  ����t�M�PHQV�҃�^]� U��Vh�DjLhD ����  ����u^]� �M�PLQV�҃�^]� �����������U��Vh�DjPhD ���y�  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�DjThD ���<�  ����u^Ë@TV�Ѓ�^���������U��Vh�DjXhD ���	�  ����t�M�PXQV�҃�^]� U��Vh�Dh�   hD �����  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�Dh�   hD ����  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�Dh�   hD ���6�  ����u^]� �M���   QV�҃�^]� �����U��Vh�Dh�   hD �����  ����u^]� �M���   QV�҃�^]� �����U��Vh�Dh�   hD ����  ����u^]� �M���   QV�҃�^]� �����U��Vh�Dh�   hD ���v�  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�Dh�   hD �5�  ����u��D�H�u�Q`V�҃���^��]ËM���   WQ�U�R�Ћ�D�Q�u���B`V�Ћ�D�Q�BpVW�Ћ�D�Q�Jl�E�P�у�_��^��]��U��Vh�Dh�   hD ��覿  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�Dh�   hD ���V�  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�Dh�   hD ����  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�Dh�   hD ���־  ����t���   ��t�MQ����^]� 3�^]� �Vh�Dh�   hD ��虾  ����t���   ��t��^��3�^����������������U��Vh�Dh�   hD ���V�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�Dh�   hD ����  ����t���   ��t�MQ����^]� ��������U��Vh�Dh�   hD ���ƽ  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������VW��3����$    �h�DjphD �o�  ����t�@p��t	VW�Ѓ����D�8 tF��_��^�������U��SW��3�V��    h�DjphD ��  ����t�@p��t	WS�Ѓ����D�8 tkh�DjphD ��  ����t�@p��tWS�Ѓ������Dh�DjphD 込  ����t�@p��t�MWQ�Ѓ����D�;uG�c����E^��t�8��~=h�DjphD �t�  ����t�@p��t	WS�Ѓ����D�8 u_�   []� _3�[]� U��Vh�Dj\hD ���)�  ����t3�@\��t,V��h�DjxhD ��  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�Dj\hD ���ɻ  ����t3�@\��t,V��h�DjdhD 觻  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�Dj\hD ���f�  ����tG�@\��t@V�ЋEh�DjdhD �E��E�    �E�    �0�  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�Dj\hD ����  ����t\�@\��tUV��h�DjdhD �Ǻ  ����t�@d��t
�MQV�Ѓ�h�DjhhD 螺  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�Dj\hD ���Y�  ������   �@\��t~V��h�DjdhD �3�  ����t�@d��t
�MQV�Ѓ�h�DjhhD �
�  ����t�@h��t
�URV�Ѓ�h�DjhhD ��  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�DjthD ��覹  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�Dj`hD �n�  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh�D���_�����^��]� ������U���Vh�Dh�   hD ����  ����tR���   ��tH�MQ�U�R���ЋuP������h�Dj`hD �ڸ  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t��D���   P�B@��]� �E��t��D���   P�BD��]� ��D���   R�PD��]� �����U�졨D�P@���   ]��������������U�졨D�P@���   ]��������������U�졨D�P@���   ]��������������U�졨D�P@���   ]��������������U�졨D���   ���   ]�����������U�졨D���   ���   ]����������̡�D�P@���   �ࡨD�P@���   ��U�졨D�P@���   ]�������������̡�D�P@���   �ࡨD���   �Bt��U�졨D�P@���   ]�������������̡�D�P@���   ��U�졨D�P@���   ]��������������U�졨DV��H@�Q$V�ҋM����t��#�����D�Q@P�B V�Ѓ�^]� �̡�D�PH���   Q�Ѓ�������������U�졨D�P@�EPQ���   �у�]� ̡�D�P@���   Q�Ѓ������������̡�D�P@�B,Q�Ѓ����������������U�졨D�P@�EPQ�J(�у�]� ����U�졨D�P@�EP�EP�EPQ�JP�у�]� ������������U�졨D�P@�EPQ�JT�у�]� ����U�졨D�P@�EP�EPQ�JX�у�]� U�졨D�P@�EPQ�J\�у�]� ����U�졨D���   �R]��������������U�졨D���   �R]��������������U�졨D���   �R ]��������������U�졨D���   ���   ]�����������U�졨D�E���   �E���   P�EP�EQ�$P�EP�EP��]� �����������U�졨D���   ���   ]����������̡�D���   �B$�ࡨD�H@�Ql�����U�졨D�H@�Apj�URj �Ѓ�]����U�졨D�H@�Apj�URh   @�Ѓ�]�U�졨D�H@�U�E�IpRPj �у�]�̡�D���   ����U��V�u���t��D���   P�B�Ѓ��    ^]�����̡�D���   �Q ��U��V�u���t��D���   P�B(�Ѓ��    ^]�����̡�D�H@�Ql�����U��V�u���t��D�Q@P�BH�Ѓ��    ^]���������U�졨D�H@���   ]��������������U��V�u���t��D�Q@P�BH�Ѓ��    ^]��������̡�D�PH���   Q�Ѓ�������������U�졨D�PH�EPQ���  �у�]� �U�졨D�H �Id]�����������������U��}qF u?V�u��t6��D���   �BDW�}W���ЋM��D�B@VQ�HhW�у����s  _^]���̡�D�P@���   ��U�졨D�P@���   ]��������������U�졨D�P@���   ]�������������̡�D�P@���   ��U�졨D���   ���   ]�����������U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U�졨D�PL�E��L  PQ�MQ�҃�]� ������������̡�D�PD�BQ�Ѓ���������������̡�D�PD�BQ�Ѓ���������������̡�D�PD�BPQ�Ѓ���������������̡�D�PD�BQ�Ѓ���������������̡�D�PD�B(Q�Ѓ����������������U�졨D�PX��Q�
�E�P�ы�M��P�@�Q�A������]� �����������U�졨D�PX��Q�J�E�P�ы�M��P�@�Q�A������]� ����������U�졨D�PX��Q�J�E�P�ы�M��P�@�Q�A������]� ����������U�졨D�PX��0VWQ�J�E�P�ы��E���   ���_^��]� �������������U�졨D�PX��0VWQ�J�E�P�ы��E���   ���_^��]� �������������U�졨D�PX�EPQ�J�у�]� ����U�졨D�PX�EPQ�J�у�]� ����U�졨D�PX�EPQ�J�у�]� ����U�졨D�PX�EPQ�J �у�]� ����U�졨D�PX�EPQ�J8�у�]� ����U�졨D�PX�EPQ�J(�у�]� ����U�졨D�PD�EP�EPQ�J,�у�]� U�졨D�HD�U�j j R�Ѓ�]�����U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U�졨D�HD�U�j j R�Ѓ�]�����U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U�졨D�U�HD�E�	Rj P�у�]���U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U�졨D�HD�U�j j R�Ѓ�]�����U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U��U��D�HD�Rj h'  �Ѓ�]��U�졨D�H@�AHV�u�R�Ѓ��    ^]�������������̡�D�HD�j j h�  �҃���������U�졨D�H@�AHV�u�R�Ѓ��    ^]�������������̡�D�HD�j j h:  �҃���������U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U���3��E��E���D���   �R�E�Pj�����#E���]�̡�D�HD�j j h�F �҃���������U�졨D�H@�AHV�u�R�Ѓ��    ^]�������������̡�D�HD�j j h�_ �҃���������U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U��E����u��]� �E���D�E�    ���   �R�E�Pj������؋�]� ̡�D�PD�BLQ�Ѓ����������������U��U��t�M��t�E��tPRQ�p�  ��]������������U�졨D�E�PH�B Q�$Q�Ѓ�]� �U�졨D�PH�EPQ���   �у�]� �U�졨D�PH��0VWQ�JP�E�P�ы��E���   ���_^��]� �������������U�졨D�PH��0VWQ�JT�E�P�ы��E���   ���_^��]� �������������U�졨D�PH�EPQ���  �у�]� �U�졨D�PH�EPQ��   �у�]� �U�졨D�PH�EP�EPQ��D  �у�]� �������������U�졨D�PH�EP�EPQ��H  �у�]� ������������̡�D�PH���  Q�Ѓ�������������U�졨D�PH�EPQ���  �у�]� ̡�D�PH�Bdj Q�Ѓ��������������U�졨D�PH�EPj Q�Jh�у�]� �̡�D�PH�BdjQ�Ѓ��������������U�졨D�PH�EPjQ�Jh�у�]� �̡�D�PH�BdjQ�Ѓ�������������U�졨D�PH�EPjQ�Jh�у�]� ��U�졨D�PH�EP�EPQ���   �у�]� �������������U�졨D�PH�EP�EPQ���   �у�]� ������������̡�D�PH�BtQ�Ѓ����������������U�졨D�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���P���������t�E��D�QH���   PVW�у���_^]� �����U��EVW���MPQ����������t�M��D�BH���   QVW�҃���_^]� ̡�D�PH��  Q�Ѓ������������̡�D�PH��  Q�Ѓ�������������U�졨D�PH�EPQ��  �у�]� �U�졨D�PH�EPQ��  �у�]� �U�졨D�PH�EP�EPQ��P  �у�]� �������������U�졨D�PH�EP�EPQ��  �у�]� ������������̡�D�PH���  Q�Ѓ������������̡�D�PH���  Q�Ѓ������������̡�D�PH���  Q�Ѓ������������̡�D�PH��   Q�Ѓ������������̡�D�PH��$  Q�Ѓ�������������U�졨D�PH�EP�EPQ��(  �у�]� �������������U�졨D�PH�EP�EP�EPQ��,  �у�]� ���������U�졨D�PH�EPQ��<  �у�]� ̡�D�PH��t  Q�Ѓ�������������U�졨D�PH�EP�EPQ��@  �у�]� �������������U�졨D�PH�EPQ��h  �у�]� ̡�DV��H@�QhWV�҃�j h�  ���=^  ����D�HH���   h�  V�҃���
��t_3�^Ë�_^��������������̡�D�P@�BhQ�Ѓ�j h�  ���]  �U�졨D�E�PH�E��,  ��P�EPQ�$Q�M�Q�ҋ�M��P�@�Q�A������]� ��������U�졨D�E�PH�E��0  ��P�EPQ�$Q�M�Q�ҋ�M��P�@�Q�A������]� ��������U�졨D�PH�EP�EPQ��4  �у�]� ������������̡�D�PH��8  Q��Y��������������U�졨D�E�PH��<  Q�$Q�Ѓ�]� �������������̡�D�PH��@  Q�Ѓ�������������U�졨D�PH�EP�EPQ��D  �у�]� �������������U�졨D�E�PH�EP�EQ�$PQ��H  �у�]� �����̡�D�PH���  Q�Ѓ������������̡�D�PH��L  Q�Ѓ������������̋��     �������̡�D�PH����  jP�у���������U�졨D�UV��HH���  R��3Ƀ������^��]� ��̡�D�PH����  j P�у��������̡�D�PH��h  Q�Ѓ������������̡�D�PH��l  Q�Ѓ������������̡�D�PH��p  Q�Ѓ�������������U�졨D�PH��Q��t  �E�P�ы�M��P�@�Q�A������]� ������̡�D�PH��x  Q�Ѓ�������������U�졨D�PH�EPQ��|  �у�]� �U�졨D�E�PH���  Q�$Q�Ѓ�]� ��������������U�졨D�E�PH���  Q�$Q�Ѓ�]� ��������������U�졨D�E�PH���  Q�$Q�Ѓ�]� ��������������U�졨D�PH�EPQ���  �у�]� �U�졨D�E�HH�U�ER�UP�EQ�$R�UP���   R�Ѓ�]��������������U�졨D�E�HH�U�ER�UQ���   �$P�ERP�у�]��U���E�M�@���  �M;�|�M;�~��]�����������U�졨D�HH�U�ER�UP���   R�Ѓ�]������������̡�D�PH���   Q��Y�������������̡�D�PH���   Q�Ѓ������������̡�D�PH���   Q��Y��������������U�졨D�PH�EP�EPQ���   �у�]� �������������U�졨D�PH�EP�EP�EP�EP�EPQ���  �у�]� ̋�� L�@    ��L��D�Px�A�JP��Y��������U�졨DV��Hx�V�AR�ЋE����u
�   ^]� ��D�Qx�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË�D�QxP�B�Ѓ�������U�졨D�Px�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U�졨D�E�HH�U�ER�UQ�$P���  R�Ѓ�]������U�졨D�HH���  ]��������������U�졨D�HH���  ]��������������U�졨D�E(�HH�U,�E$R�U Q�$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�(]��������������U�졨D�HH���  ]��������������U�졨D�E�PH�EPQ�$Q���  �у�]� ����������U���SV����  �؉]����   �} ��   ��D�HH���  j h�  V�҃��E��u
^��[��]� �MW3��}�� �  ����   �]��I �E�P�M�Q�MW�ߝ  ��ta�u�;u�Y�I ������u�E�������L�;Ht-��D�Bx�S�@����QR�ЋD������t	�M�P�Ü  F;u�~��}��MG�}�莜  ;��v����]�_^��[��]� ^3�[��]� ��������������U�����DSV�ًHH���  j h�  S�]��ҋ�����u
^3�[��]� �E��u��D�HH���  �'��u��D�HH���  ���uš�D�HH���  S�ҋȃ��E��t�W褛  ��D�HH���   h�  S3��҃����  ���_�u����    ��D�Hx�U�B�IWP�ы�������   ��D�F�J\�UP�A0R�Ѓ���t�K�Q�M�u�  ��D�F�J\�UP�A0R�Ѓ���t�K�Q�M�L�  �E��;Pt&�F��D�Q\�J0P�EP�у���t	�MS��  ��D�v�B\�M�P0VQ�҃���t�M�CP��  ��D�QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U�졨D�HH��  ]�������������̡�D�PH��  Q��Y��������������U�졨D�HH���  ]��������������U��Q��V�uW�}Q�$V���T  �]��E��E������Au������E������{����]Q�E���$V�X  _^��]���������U��� ��V�u�U�W�U��}�]�E�PV�M�Q����S  �E��E�����E��Au���U��������z�����U����E�������z���U�����]���������Au@�����U����E�������z0�����]�U��ER�]�V�E����]��E��]���W  _^��]��]�����������Au����������U�졨D�HH�U�j R�Ѓ�]�������U�졨D�H@�AHV�u�R�Ѓ��    ^]�������������̡�D�HH�j h�  �҃�����������U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U�졨D�HH�Vj h  �ҋ�������   �EPh�  ��������t]��D�QHj P���   V�ЋMQh(  ��������t3��D�JH���   j PV�ҡ�D���   �B��j j���Ћ�^]á�D�H@�QHV�҃�3�^]�����U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U�졨D�HH�Vj h�  �ҋ�����u^]á�D�HH�U�E��(  RPV�у���u��D�B@�HHV�у�3���^]�����U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U�졨D�HH�I]�����������������U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U�졨D�PH�EPQ���  �у�]� �U�졨D�PH�EPQ���  �у�]� ̡�D�PH���  Q�Ѓ�������������U�졨D�HH���  ]��������������U�졨D�E�HH�U(�E$R�U P�ER�UP�ER�U���\$�E�$P��p  R�Ѓ�$]������������̡�D�PH��  Q�Ѓ�������������U�졨D�PH�EP�EPQ��  �у�]� ������������̡�D�PH��8  Q�Ѓ�������������U�졨D�PH�EP�EP�EPQ��   �у�]� ��������̡�D�PH��$  Q�Ѓ������������̡�D�PH��(  Q�Ѓ�������������U�졨D�PH�EPQ��0  �у�]� �U�졨D�PH�EPQ��4  �у�]� ̋������������������������������̡�D�HH��  ��U�졨D�HH��  ]��������������U�졨D�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��  �у�0]�, ���������U�졨D�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��x  �у�0]�, ���������U�졨D�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��  �у�0]�, ���������U�졨D�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��|  �у�0]�, ��������̡�D�PH��X  Q�Ѓ�������������U�졨D�PH�EPQ���  �у�]� ̡�D�PH���  Q�Ѓ�������������U�졨D�HH��\  ]��������������U�졨D�HH��d  ]��������������U�졨D��W���HH���   j h�  W�҃��} u�   _��]� Vh�  ����������tq��D�HH���   j VW�҃��M��G  �EPh�  �M���O  �EQ�$h�  �M��"P  ��D�Q@�Jdj �E�PV�у��M���G  ^�   _��]� ^3�_��]� �����������U��S�]�; VW��u7��D�U�HH���   RW�Ѓ���u��D�QH���   jW�Ѓ���t�   �����   ��D�QH���   W�Ѓ��} u(��D�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;��D�U�HH�ER�USP���  VRW�Ћ�D���   �B(�����Ћ���uŃ; u��D�QH���   W�Ѓ���t3���   �W��u1��D�QH���   �Ћ�D�E�QH���   PW�у�_^[]� ��D�BH���   �у��} u0��D�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ��D�QH�j h  �Ћ؃���u_^[]� ��D���   �u�Bx���Ћ�D���   P�B|���Ѕ�t_���$    ���D�E�QH�MP�Ej Q���  VPW�у���t��D���   �ȋBHS�Ћ�D���   �B(���Ћ���u�_^��[]� ��U��EV���u��D�HH���  �'��u��D�HH���  ���u��D�HH���  V�҃���u3�^]� P�EP������^]� ���������U���@��D�HH���   SV�uWh�  V�ҋ���D�HH�Q|3�Sh�  V�}��]��҉E�3����E�E��E�;���  ��D���   �B���Ћ�D=�  �  �QH�Bx3�Wh:  V�Ћ�D�QH�E䋂�   h�  V�Ћ�D�QHW�؋B|h�  V�]ԉ}��Ћ�D�QH�E苂8  V�Ћ�D�QH�EЋ�$  V�Ѓ�(�E��E�X��~{�M���M܋MЅ�tMj�W�Y�  ���t@�@�Ẽ|� ��~����%�������;�u/���ر  ;E�~�E؋�虱  E���E܋;Pu�E���E��E�G;}�|��}� tm�}�j V���3�������   ���������tM���y����]�;�uB��D�H��H  �<[j ��j W�҃��E����   �M�WP�~���P�X�������]ࡨD�H��H  �<[3�S��SW�҃��E�;�tr�M�;�t;�tWQP觺  ���E�;�~!��D�QS��SP��H  �Ѓ��E�;�t4��D�E��QH��(  j�PV�у���t�}�;�tAjV���<�����u'�U�R��p  �E�P��p  �M�Q��p  ��_^3�[��]Ë�������E���]���D�BH�H|Sh�  V�у�3�9]ԉE�]���  �}���I �MЅ��  j�S�m�  �����  �@�Ẽ|� ���U�~�
���%�������;��  3�3�9J�M���   �����������tz�]��U���������M���ʋ���]��U��҉T��]�@�U؋Q�T��]��U�@B�T��Q�]�@�T��U؋]�@���T��I�U�@�L��M؋U�@@�����U�@�M�A;J�M��e����E܅��h  �+�j��P�E�P�M���  �M�v���E��E�3�+��E����    �}� �M����E�t-�M�@���MĉU؋U�ʋU؋��U؋R�Q�U؋R�Q;]܋U��@����M؋M���U؋R�Q�U؋R�Q}j����    �E��M�9�uU�ыL�����������w4�$�<� �M����4�"�U����t��M����t�
�U����t��;]�|��E�F;]��"����S  ��M�3�;G�Å���   �E��v���W��R�����Q�P�I�H�O��I�M����P�Q���P�I�H��@�E���U��Lv�����P�Q�@�A��t&�G�U�@���U��Lv	�����P�Q�@�A�G��U��@���U�v�����P�Q�@�A�G��w��U��@���U�F�v�����P�Q�@�A��w��U�F�@���U�v�����P�Q�@�A�7F��t+�G�U��@���U�v�����P�Q�@�A�wF���O�]�C��;]ԉ]�������U�R��l  �E�P��l  ���  ���   �B����=  ��  ��D�QH�B|j h(  V�Ћ�D�QH�����   h(  V�ЋЃ�3��U؅�~�ǅ�t�|� t�K��\K�@;�|�]��]���D�Q��H  �[j ��j S�Ѓ��E�����   �}� t��t�M�SQP薵  ���]؋�D�B��H  �j ��j S�у��E��tP��t��tSWP�Z�  ���M����+�D�RH��PQ�E���  V�Ѓ���u�M�Q��k  �U�R�k  ��_^3�[��]á�D�HH�Q|j h�  V�҉E���D�HH�Q|j h(  V��3�3�3ۃ�9U؉Eĉ}̉]���   �u荛    �ޅ���   ���E�    ~g�u�<�R��   ����d$ �u��>��\>��EԉY�v�q�u��\7�t7�Y�^���Y�v�]�q�u�B@B����;�|��}̃|� tO�Eԋu�8�E��I���R�4����A�F�I�N�M��u���B�R�4����A�F�I�N�u�B<މ}�C;]؉]������M�3�3�;�~�Uĉt���   @;�|�U�R�Rj  ���E�P�Fj  ��_^�   [��]ÍI �{ �{ �{ �{ ����U��E� �M+]� ���������������U��V��V�L��D�Hx�AR�Ѓ��Et	V�n  ����^]� ���������̡�D�H8�������U�졨D�H8�AV�u�R�Ѓ��    ^]��������������U�졨D�P8�EP�EPQ�J�у�]� U�졨D�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U�졨D�P8�EP�EPQ�J�у�]� U�졨D�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H�A0]�����������������U�졨D�H�I4]�����������������U�졨D�H�Q`V�uV�ҡ�D�H�Q<V�҃���^]�����̡�D�H�Q@�����U�졨D�H�ID]����������������̡�D�H�QH����̡�D�H�QL�����U�졨D�H�AP]�����������������U�졨D�H�AT]�����������������U�졨D�H���  ]��������������U�졨D�H��|  ]��������������U�졨D�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡�D�H���   �⡨D�H��   ��U�졨D�H�U�ER�UP�ER�UP���   Rh�*  �Ѓ�]����������������U�졨D�H�A]�����������������U�졨D�H�Ad]�����������������U�졨D�H�Ah]�����������������U�졨D�H�Al]����������������̡�D�H�Qp����̡�D�H�Qt����̡�D�H�Qx�����U�졨D�H�A|]�����������������U�졨D�H���   ]��������������U�졨D�H���   ]��������������U�졨D�H���  ]��������������U�졨D�H��X  ]��������������U�졨D�H���   ]��������������U�졨D�H���  ]��������������U��V�u���B  ��D�H�U���   VR�Ѓ���^]������U�졨D�H���   ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]�������������̡�D�H���   ��U�졨D�H���  ]��������������U�졨D�H��P  ]��������������U�졨D�H��T  ]��������������U��V�u���4  ��D�H���   V�҃���^]���������̡�D�H���  ��U�졨D�H��\  ]��������������U�졨D�H�U���   ��R�E�P�ы�M��P�@�Q�A������]�������U�졨D�H��  ]��������������U��U�E��D�H�E���   R���\$�E�$P�у�]�U�졨D�H���   ]��������������U�졨D�H��   ]��������������U�졨D�H��h  ]��������������U�졨D�H��l  ]��������������U�졨D�H��  ]��������������U�졨D�H���  ]��������������U�졨D�H��$  ]��������������U�졨D�H��(  ]��������������U�졨D�H��,  ]��������������U�졨D�H��0  ]��������������U�졨D�H��4  ]��������������U�졨D�H��8  ]��������������U�졨D�H��<  ]��������������U�졨D�H��@  ]��������������U�졨D�P���E�P�E�P�E�PQ��D  �у����#E���]����������������U�졨D�P���E�P�E�P�E�PQ��D  �у����#E���]����������������U�졨D�P���E�P�E�P�E�PQ��D  �у����#E���]����������������U�졨D�H���  ]��������������U��V�u(V�u$�E�@��D�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@��D�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U�졨D�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�졨D�P0�EP�EP�EP�EPQ���   �у�]� ����̡�D�P0���   Q�Ѓ�������������U�졨D�P0�EP�EPQ���   �у�]� �������������U�졨D�P0�EP�EP�EP�EPQ���   �у�]� ����̡�D�P0���   Q�Ѓ������������̡�D�H0���   ��U�졨D�H0���   V�u�R�Ѓ��    ^]�����������U�졨D�H���  ]��������������U�졨D�H���  ]�������������̡�D�H���  �⡨D�H��  ��U�졨D�H��,  ]��������������U�졨D�H��8  ]��������������U�졨D�H��0  ]��������������U�졨D�H��(  ]��������������U�졨D�H��H  ]��������������U�졨D�H�U�E���  ��VR�UPR�E�P�ыu�    �F    ��D���   �Qj PV�ҡ�D���   ��U�R�Ѓ� ��^��]��������U���Vj hLGOg�M���-  P�E�hicMCP�k������M��0.  ��D���   �JT�E�P�у���u(�u���z-  ��D���   ��M�Q�҃���^��]á�D���   �AT�U�R�Ћu��P���-  ��D���   �
�E�P�у���^��]�������������U�졨D�H��`  ]��������������U�졨D�H���  ]��������������U�졨D�H�U���  ��V�uVR�E�P�у����  �M��  ��^��]�����U�졨D�H���  ]��������������U�졨D�H�U���  ��VWR�E�P�ы�D�u���B�H`V�ы�D�B�HpVW�ы�D�B�Pl�M�Q�҃�_��^��]����������������U�졨D�H�U���  ��VWR�E�P�ы�D�u���B�H`V�ы�D�B�HpVW�ы�D�B�Pl�M�Q�҃�_��^��]����������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H��   ]��������������U�졨D�H��  ]��������������U�졨D�H��  ]��������������U��E�M�U��VWPQR�����     �@    ��D���   �M�Rj QP�ҡ�D�H���  �U���R�Ћ�D�Q�u���B`V�Ћ�D�Q�BpVW�Ћ�D�Q�Jl�E�P�у�(_��^��]�����������U�졨D�H�U�E��  ��VR�UPR�E�P�ыu�    �F    ��D���   �Qj PV�ҡ�D���   ��U�R�Ѓ� ��^��]��������U���  �13ŉE��M�EPQ������R�Ӧ  ��D�H���  ������Rh\�ЋM�3̓�肟  ��]�������������U�졨D�H��h  ��V�U�WR�Ћ�D�Q�u���B`V�Ћ�D�Q�BpVW�Ћ�D�Q�Jl�E�P�у�_��^��]����U�졨D�H��l  ��V�U�WR�Ћ�D�Q�u���B`V�Ћ�D�Q�BpVW�Ћ�D�Q�Jl�E�P�у�_��^��]����U�졨D�H���  ���҅�tbh���M��(  �EPh���M���0  �MQh���M���0  j �U�R�E�hicMCP�#�����D���   �
�E�P�у��M���(  ��]�U�졨D�H���  ��V�҅�u��D�H�u�Q`V�҃���^��]�Wh!���M��(  �EPh!���M��K0  j �M�Q�U�hicMCR������D���   P�BH�Ћ�D�Q�u���B`V�Ћ�D�Q�BpVW�Ћ�D���   �
�E�P�у�$�M��(  _��^��]�����������U�졨D�H���  ���҅�u��]�Vh#���M��d'  �EPh#���M��/  j �M�Q�U�hicMCR�������D���   P�B8�Ћ�D���   �
���E�P�у��M��|'  ��^��]������U�졨D�H���  ���҅�u��]�Vhs���M���&  �EPhs���M��/  j �M�Q�U�hicMCR�O�����D���   P�B8�Ћ�D���   �
���E�P�у��M���&  ��^��]������U�졨D�H��,  ]��������������U�졨D�H���  ]��������������U�졨D�H��0  ]��������������U��V�u���t��D�QP���  �Ѓ��    ^]������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]�������������̡�D�H���  ��U�졨D�H���  ]��������������U�졨D�H���  ]�������������̡�D�H���  ��U�졨D�H�U���  ��VR�E�P�ыu��P����$  �M���$  ��^��]�����U�졨D�H���  ]��������������U�졨D�H��   ]��������������U�졨D�H��  ]��������������U�졨D�H��  ]��������������U�졨D�H��  ]��������������U�졨D�H��  ]��������������U���h����M��#  j �E�P�M�hicMCQ�9�����D���   ��M�Q�҃��M���#  ��]�������U�졨D�H��   ]��������������U�졨D�H���  ]��������������U�졨D�H��L  ]�������������̡�D�H��P  ��U�졨D�H��T  ]������������������������������U�졨D�H��|  ]��������������U�졨D�H�A`�U��� R�Ћ�D�Q�Jdj j��E�h`P�ыUR�E�P�M�Q轟����D�B�Pl�M�Q�ҡ�D�H�A�U�R�Ћ�D�Q�Jl�E�P�у�,��]��U�졨D�P�EP�EP�EPQ�Jd�у�]� �����������̡�D�H$�Q�����U�졨D�H$�U�AR�Ѓ�]��������U�졨D�H$�A]����������������̡�DV��H$�QDV�҃���^���������U�졨DV��H$�QDV�ҡ�D�U�H$�AdRV�Ѓ���^]� U�졨DV��H$�QDV�ҡ�D�U�H$�ARV�Ѓ���^]� U�졨DV��H$�QDV�ҡ�D�H$�U�ALVR�Ѓ���^]� ��D�P$�BHQ��Y�U�졨D�P$�EPQ�JL�у�]� ���̡�D�P$�BQ�Ѓ����������������U�졨D�P$�EP�EP�EPQ�J�у�]� ������������U�졨D�P$�EP�EP�EPQ�J�у�]� �����������̡�D�P$�BQ�Ѓ����������������U�졨DVW�}��H�Q`W�ҡ�D�H$�QV�ҋ�����t ��D�H�QpWV�ҡ�D�H�QV�҃���_^]� ���������U�졨D�P$�EPQ�J�у�]� ���̡�D�P$�B(Q��Yá�D�P$�BhQ��Y�U�졨D�P$�EPQ�J,�у�]� ����U�졨D�P$�EPQ�J0�у�]� ����U�졨D�P$�EPQ�J4�у�]� ����U�졨D�P$�EPQ�J8�у�]� ����U�졨D�UV��H$�ALVR�Ѓ���^]� ��������������U�졨D�H$�QDV�uV�ҡ�D�H$�U�ALVR�Ћ�D�E�Q$�J@PV�у���^]���������������U�졨D�UV��H$�A@RV�Ѓ���^]� ��������������U�졨D�P$�EPQ�J<�у�]� ����U�졨D�P$�EPQ�J<�у����@]� ���������������U��V�u���t��D�Q$P�B�Ѓ��    ^]���������U�졨D�P$�EP�EPQ�JP�у�]� U�졨D�P$�EPQ�JT�у�]� ���̡�D�H$�QX�����U�졨D�H$�A\]�����������������U�졨D�P$�EP�EP�EPQ�J`�у�]� �����������̡�D�H(�������U�졨D�H(�AV�u�R�Ѓ��    ^]��������������U�졨D�P(�EP�EP�EP�EP�EP�EPQ�J�у�]� ��D�P(�BQ�Ѓ����������������U�졨D�P(�EPQ�J�у�]� ����U�졨D�P(�EP�EP�EPQ�J�у�]� ������������U�졨D�P(�EP�EPQ�J�у�]� U�졨D�P(�EjP�EPQ�J�у�]� ��������������U�졨D�P(�EP�EPQ�J�у�]� ��D�P(�B Q�Ѓ���������������̡�D�P(�B$Q�Ѓ���������������̡�D�P(�B(Q�Ѓ����������������U�졨D�P(�EPQ�J,�у�]� ����U�졨D�P(�EPQ�JP�у�]� ����U�졨D�P(�EPQ�JT�у�]� ����U�졨D�P(�EPQ�JX�у�]� ����U�졨D�P(�EPQ�J\�у�]� ����U�졨D�P(�EPQ�J`�у�]� ����U�졨D�P(�EPQ�Jp�у�]� ����U�졨D�P(�EPQ�Jd�у�]� ����U�졨D�P(�EPQ�Jh�у�]� ����U�졨D�P(�EPQ�Jl�у�]� ����U�����DV���E�    �E�    �H(�A`�U�RV�Ѓ�����   �E���uI��D�Q�J`�E�P�ы�D�B�M�@pQ�U�R�Ћ�D�Q�Jl�E�P�у��   ^��]� ��D�J��H  j j P�҃��E���u��D�H(�Q,j�V�҃�3�^��]� ��D�Q(�M��Rj QPV�҃���u�E�P�:H  ��3�^��]� �M��U�j IQ�MR�����E�P�H  ���   ^��]� ���U�졨D��V��H�A`�U�R�Ѓ��M�Q������^��u��D�B�Pl�M�Q�҃�3���]� ��D�H$�E�I�U�RP�ы�D�B�Pl�M�Q�҃��   ��]� �U��Q��D�P(�E�PQ�JP�у���u��]� �E3�8U���   ��]� �����U�졨DVW�}��H(�QhWV�҃���t$��D�H(�Qh��WV�҃���t_�   ^]� _3�^]� ����U�졨DVW�}��H(�QhWV�҃���t>��D�H(�Ah�WRV�Ѓ���t%��D�Q(�Bh��WV�Ѓ���t_�   ^]� _3�^]� ����������U�졨DVW�}��H(�QlWV�҃���t>��D�H(�Al�WRV�Ѓ���t%��D�Q(�Bl��WV�Ѓ���t_�   ^]� _3�^]� ����������U��VW�}W��������t8�GP��������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U�졨D�P(�EPQ�J0�у�]� ����U�졨D�P(�EPQ�J4�у�]� ����U�졨D�P(�EPQ�J8�у�]� ����U�졨D�P(�EPQ�J<�у�]� ����U�졨D�P(�EPQ�J@�у�]� ����U�졨D�P(�EP�EPQ�Jt�у�]� U�졨D�P(�EPQ�JD�у�]� ����U�졨D�E�P(�BHQ�$Q�Ѓ�]� �U�졨D�E�P(�BL���$Q�Ѓ�]� ��������������̡�D�H,�Q����̡�D�P,�B8�����U�졨D�H,�A V�u�R�Ѓ��    ^]�������������̡�D�P,�B<�����U�졨D�P,�R@��VW�E�P�ҋu����D�H$�QDV�ҡ�D�H$�QLVW�ҡ�D�H$�AH�U�R�Ѓ�_��^��]� �������U�졨D�P,�E�RH��VWP�E�P�ҋu����D�H�Q`V�ҡ�D�H�QpVW�ҡ�D�H�Al�U�R�Ѓ�_��^��]� ��̡�D�H,�j j �҃��������������U�졨D�P,�EP�EPQ�J�у�]� U�졨D�H,�AV�u�R�Ѓ��    ^]�������������̡�D�P,�BQ�Ѓ���������������̡�D�P,�BQ�Ѓ���������������̡�D�P,�BQ�Ѓ���������������̡�D�P,�B,����̡�D�P,�BD����̡�D�P,�B0�����U�졨D�P,�R4]�����������������U�졨D�H,�A$]�����������������U�졨D�H,�AL]�����������������U�졨D�H,�A(]�����������������U�졨DVW�}��H$�QDW�ҡ�D�H,�QV�ҋ�����t ��D�H$�QLWV�ҡ�D�H$�QV�҃���_^]� ���������U�졨D�H�I]�����������������U�졨D�H�A]�����������������U�졨D�H�I]�����������������U�졨D�H�A]�����������������U�졨D�H�I]�����������������U�졨D�H��\  ]��������������U�졨D�H�A ]�����������������U�졨D�H�A$]�����������������U�졨D�H�I,]�����������������U�졨D�H��p  ]��������������U�졨D�H��t  ]��������������U�졨D�H��x  ]��������������U�졨D�H$�QDVW�}W�ҡ�D�H�Q(���ҋ���t ��D�H$�QLWV�ҡ�D�H$�QV�҃���_^]���������������U�졨D�H$�QDVW�}W�ҡ�D�H��X  ���ҋ���t ��D�H$�QLWV�ҡ�D�H$�QV�҃���_^]������������U�졨D�H��d  ]��������������U�졨D�H�U��L  ��VWR�E�P�ы�D�u���B$�HDV�ы�D�B$�HLVW�ы�D�B$�PH�M�Q�҃�_��^��]����������������U��V�ujV��������^]���������̡�D�H���   ��U�졨D�H���   V�uV�҃��    ^]�������������U�졨D�P�EP�EP�EPQ���   �у�]� ��������̡�D�P���   Q�Ѓ������������̡�D�P���   Q�Ѓ�������������U�졨D�P�EPQ�JL�у�]� ����U�졨D�P�EPQ�JP�у�]� ����U�졨D�P�EPQ�JT�у�]� ����U�졨D�P�EPQ�JX�у�]� ����U�졨D�P�EPQ�J\�у�]� ����U�졨D�P�EPQ�J`�у�]� ����U�졨D�P�EPQ���   �у�]� �U�졨D�P�EPQ�Jd�у�]� ����U�졨D�P�EPQ�Jh�у�]� ����U�졨D�P�EPQ�Jl�у�]� ����U�졨D�P�EPQ�Jp�у�]� ����U�졨D�P�EPQ�Jt�у�]� ����U�졨D�P�EPQ�Jx�у�]� ����U�졨D�P�EPQ�J|�у�]� ����U�졨D�P�EPQ���   �у�]� �U�졨D�P�EPQ���   �у�]� �U�졨D�P�EPQ���   �у�]� �U�졨D�P�EPQ���   �у�]� �U�졨D�P�EP�EPQ���   �у�]� �������������U�졨D�P�EP�EPQ���   �у�]� �������������U�졨D�P�EPQ���   �у�]� �U��E��t ��D�R P�B(Q�Ѓ���t	�   ]� 3�]� U�졨D�P �E�RhQ�MPQ�҃�]� U��E��u]� ��D�R P�B,Q�Ѓ��   ]� ������U�졨D�P�EPQ�
�у�]� �����U�졨D�P�EPQ�J�у�]� ����U�졨D�P�EPQ�J�у�]� ����U�졨D�P�EPQ�J�у�]� ����U�졨D�P�EPQ�J�у�]� ����U�졨D�P�EPQ�J�у�]� ����U�졨D�P�EP�EPQ���   �у�]� �������������U�졨D�E�P�BQ�$Q�Ѓ�]� �U�졨D�E�P�B���$Q�Ѓ�]� ���������������U�졨D�P�EPQ�J �у�]� ����U�졨D�P�EPQ�J$�у�]� ����U�졨D�P�EPQ�J(�у�]� ����U�졨D�P�EPQ�J,�у�]� ����U�졨D�P�EPQ�J0�у�]� ����U�졨D�P�EPQ�J4�у�]� ����U�졨D�P�EPQ�J8�у�]� ����U�졨D�P�EPQ�J<�у�]� ����U�졨D�P�EP�EP�EP�EPQ���   �у�]� �����U�졨D�P�EPQ�JD�у�]� ����U�졨D�P�EPQ���   �у�]� �U�졨D�P�EP�EPQ�JH�у�]� ��D�P���   Q�Ѓ�������������U�졨D�P�EPQ���   �у�]� �U�졨D�P�EPQ���   �у�]� �U�졨D�P�EPQ���   �у�]� �U�졨D�P�EP�EPQ���   �у�]� ������������̡�D�P���   Q�Ѓ�������������U�졨D�P�EP�EPQ���   �у�]� ������������̡�D�P���   Q�Ѓ������������̡�D�P���   Q�Ѓ������������̡�D�P���   Q�Ѓ�������������U�졨D�H���   ]��������������U�졨D�H���   ]��������������U�졨D�H�U�E��VWRP��4  �U�R�Ћ�D�Q�u���B`V�Ћ�D�Q�BpVW�Ћ�D�Q�Jl�E�P�у�_��^��]������������U�졨D�H��8  ]��������������U�졨DVW�}��H$�QDW�ҡ�D�H$�Q V�ҋ�����t ��D�H$�QLWV�ҡ�D�H$�QV�҃���_^]� ���������U�졨DVW�}��H$�QDW�ҡ�D�H$�Q$V�ҋ�����t ��D�H$�QLWV�ҡ�D�H$�QV�҃���_^]� ���������U���V�uV�E�P�������e�����D�Q$�JH�E�P�у���^��]� �������U�졨D�P(�} ����PQ�J0�у�]� �������������U�졨DVW�}���H(�]�E�QHQ�$V�҃���t-�G��D�H(�]�E�QHQ�$V�҃���t_�   ^]� _3�^]� U�졨DVW�}���H(�]�E�QHQ�$V�҃���tO�G��D�H(�]�E�QHQ�$V�҃���t-�G��D�H(�]�E�QHQ�$V�҃���t_�   ^]� _3�^]� ��������������U�졨DVW�}���H(�QL���$V�҃���tG��D�G�H(�QL���$V�҃���t)��D�G�H(�QL���$V�҃���t_�   ^]� _3�^]� ����������U��VW�}W���������t8�GP���������t)�OQ���������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W��������t8�GP��������t)�O0Q���������t��HW���������t_�   ^]� _3�^]� ������������U�졨DS�]VW���H�QPj S�ҋ�D�H��H  j Fj V�҃��E��u��D�H(�Q,j�W�҃�_^3�[]� ��D�Qj VP�BTS�Ћ�D�Q(�B@VW�Ѓ���t"��D�E�Q(�JVPW�у���t�   �3��UR�01  ��_��^[]� ����U���V�E���MP����P���#�����D�Q�Jl���E�P�у���^��]� ���U���V�u�E�P��������D�Q$�J�E�P�у���u��D�B$�PH�M�Q�҃�3�^��]á�D�H�A�U�jR�Ѓ���u�M�Q��������t���D�H�QjV�҃���u0��D�H�Q V�҃���u��D�H$�AH�U�R�Ѓ�3�^��]Ë�D�Q$�JH�E�P�у��   ^��]�������U���<��DSVW�E�    ��t�E�P�   ���������D�Q$�JD�E�P�   �у��u���D�B$�}�HDW�ы�D�B$�HLWV�у���t��D�B$�PH�M�Q����҃���t��D�H$�AH�U�R�Ѓ���_^[��]���̡�D�H�Qj��҃���������������U�졨D�H�U�AR�Ѓ�]��������U�졨D�H�A]����������������̡�DV��H���   j�V�҃���^����U�졨D�UV��H���   RV�Ѓ���^]� �����������U�졨DV��H���   j�V�ҡ�D�H�U���   j VR�Ѓ���^]� �����̡�D�P�BQ��Y�U�졨D�UV��H���   j VR�Ѓ���^]� ���������U�졨D�P�EP�EPQ���   �у�]� �������������U�졨D�P�EP�EP�EPQ���   �у�]� ���������U�졨DVW���H�Qj��ҋ�����u_^]� �U��D�H���   RVW�Ѓ�_��^]� ����������U�졨D�P�EPQ�J�у�]� ����U�졨D�P�EPQ�J�у����@]� ��������������̡�D�P�BQ��Yá�D�P�BQ�Ѓ����������������U�졨D�P�EPQ�J�у�]� ����U�졨D�P�EPQ�Jh�у�]� ����U�졨D�P�EPQ�Jt�у�]� ����U�졨D�P�EPQ�Jl�у�]� ����U�졨D�P�EPQ�Jp�у�]� ����U�졨D�UV��H�AlRV�Ѓ����u3�^]� ��D�QP�B|V�Ѓ�^]� �U�졨D�P�EPQ�J|�у�]� ����U�졨DVW�}��H�QlWV�҃����u	�E_^]� ��D�H�QHWV�҃�_^]� ��������������U�졨DVW�}��H�QlWV�҃����u	�E_^]� ��D�H�QLWV�҃�_^]� ��������������U�졨DVW�}��H�QlWV�҃����u�E�U_^]� ��D�H���   WV�҃�_^]� ��������U�졨DVW�}��H�QlWV�҃����tI��D�H���   WV�ҋ�D���   �QV�҃���u��D���   �Q`jV�҃�_^]� �E_^]� �������������U�졨DVW�}��H�QlWV�҃����u	�E_^]� ��D�H�QDWV�҃�_^]� ��������������U�졨D��VW�}��H�QlWV�҃����u�M��E��Q�I_�P�H^��]� ��D�B�P`W�M�VQ�ҋ�M��P�@���Q_�A��^��]� ����������U�졨D��0VW�}��H�QlWV�҃����u�E�u�   ���_^��]� ��D�H�AdW�U�VR�Ћ��E���   ���_^��]� ���������U�졨D��VW�}��H�QlWV�҃����u0��D�H�u�Q`V�ҡ�D�H�U�ApVR�Ѓ�_��^��]� ��D�Q�BPWV�Ћ�D�Q�J`���E�P�у���t$��D�B�Pp�M�QV�ҡ�D�H�QV�҃���D�H�u�Q`V�ҡ�D�H�Ap�U�VR�Ћ�D�Q�Jl�E�P�у�_��^��]� �����������U�졨D��VW�}��H�QlWV�҃����u�E�uP������_��^��]� ��D�Q�BTWV�Ѓ��M�E�v����E��t	P�M������MQ������u���U�R��������M������_��^��]� ����������U�졨D�P�EVWPQ�J\�ы�D�u�����B���   j�V�х�t ��D�B���   j VW�у�_��^]� ��_��^]� ��������������U�졨D�P�EPQ�J\�у�]� ����U�졨D��VW�}��H�QlWV�҃����u�M��E�I_��H^��]� ��D�B�PXW�M�VQ�ҋ�M�@��_�A���^��]� ������U�졨D�P�EP�EPQ�J$�у�]� U�졨D�P�EP�EPQ�J(�у�]� U�졨D�P�EP�EP�EPQ���   �у�]� ���������U�졨D�E�P�EQ�$PQ�J �у�]� �������������U����E��D�E�   �E��B���   �U�R�URQ�Ћ�D���   �
�E�P�у���]� ������U�졨D�P�EP�EPQ�J<�у�]� U�졨D�P�EP�EPQ�J@�у�]� U�졨D�P�EP�EPQ�J,�у�]� U�졨D�P�EP�EPQ�J0�у�]� U�졨D�P�EP�EPQ�J8�у�]� U�졨D�P�EP�EPQ�J4�у�]� U�졨D�P�EPQ���   �у�]� �U�졨D�P�EP�EPQ���   �у�]� �������������U�졨D�P�EP�EP�EPQ���   �у�]� ���������U�졨D�P�EP�EPQ���   �у�]� �������������U�졨D�P�EPQ���   �у�]� �U�졨D�P�EPQ���   �ы�D���   �QXP�҃�]� ���������������U�졨D�P�EPQ���   �ыU�M��RQ���fi  ]� ��U�졨D�P�EP�EP�EPQ���   �у�]� ���������U�졨D�P�EP�EPQ���   �у�]� �������������U�졨D�P�Eh#  P�EPQ���   �у�]� ��������U�졨D�P�EhF  P�EPQ���   �у�]� ��������U�졨D�P�EPQ���   �ы�D���   �URP�A`�Ѓ�]� �����������U�졨D�P�EPQ���   �у�]� �U�졨D�P�EP�EPQ���   �у�]� �������������U�졨D�P�EP�EPQ���   �у�]� ������������̡�D�P���   Q��Y�������������̡�D�HL��8  ��U�졨D�H@�AHV�u�R�Ѓ��    ^]�������������̡�D�HL�������U�졨D�H@�AHV�u�R�Ѓ��    ^]�������������̡�D�PL���   Q�Ѓ�������������U�졨D�PL�EP�EPQ���   �у�]� �������������U�졨DV��HL���   V�҃���u��D�U�HL���   j RV�Ѓ�^]� ��D���   �ȋBP�Ћ�D���   �MP�BH��^]� �����̡�D�PL��p  Q�Ѓ�������������U�졨D�PL�EP�EPQ��t  �у�]� ������������̡�D�HL�Q�����U�졨D�H@�AHV�u�R�Ѓ��    ^]��������������U��V�uW�����O�����D�U�HL�AVRW�Ѓ�_��^]� �U�졨D�PL�EPQ��   �у�]� �U�졨D�PL�EP�EPQ�J�у�]� ��D�PL�B Q�Ѓ���������������̡�D�PL�B$Q�Ѓ���������������̡�D�PL�B(Q�Ѓ����������������U�졨D�PL�EP�EPQ�J,�у�]� U�졨D�PL�EPQ��|  �у�]� �U�졨D�PL�EP�EP�EPQ�J0�у�]� ������������U�졨D�PL�EP�EP�EP�EPQ�J4�у�]� �������̡�D�PL�B8Q�Ѓ���������������̡�D�PL�B<Q�Ѓ����������������U�졨D�PL�EP�EPQ��`  �у�]� ������������̡�D�PL���   Q�Ѓ�������������U�졨D�PL��VQ��   �E�P�ыu��P�������M�������^��]� �����U�졨D�PL�E��T  ��VPQ�M�Q�ҋu��P���B����M��z�����^��]� ̡�D�PL�B@Q�Ѓ���������������̡�D�PL�BDj Q�Ѓ��������������U�졨D�PL���   ]��������������U�졨D�PL���   ]��������������U�졨D�PL��4  ]��������������U�졨D�PL���   ]��������������U�졨D�PL���   ]��������������U�졨D�PL��  ]��������������U�졨D�PL���   ]��������������U�졨D�PL���   ]��������������U�졨D�PL��0  ]��������������U�졨D�PL�EPQ�JT�у�]� ���̡�D�PL�BQ��Y�U�졨D�PL�EP�EPQ�JX�у�]� U�졨D�PL�Ej PQ�J\�у�]� ��U�졨D�PL�Ej PQ�J`�у�]� ��U�졨D�PL�EjPQ�J\�у�]� ��U�졨D�PL�EjPQ�J`�у�]� ��U���SVW3��E��P�M��}��}��E��  �}�}��dz��W�M�Q�U�R���4������M����m����t��D���   ��U�R�Ѓ�_^3�[��]Ë�D���   �J8�E�P�ы�D�����   ��M�Q�҃�_��^[��]��������������U���3�V�E�E�E��P�M��E�   �E�   �E��  �y��j�M�Q�U�R��蝀���M��el����D���   ��U�R�Ѓ�^��]�����������U�����D�UVW3���}��}����   �I(R�E�P�у��U�R�M��E��  �}�}��*y��j�E�P�M�Q�������M���k����D���   ��M�Q�҃�_^��]� ��U�����D�UVW3���}��}����   �I(R�E�P�у��U�R�M��E��  �}�}��x��j�E�P�M�Q������M��ak����D���   ��M�Q�҃�_^��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��Dx��W�M�Q�U�R��������M�����j����t+�u��������D���   ��U�R�Ѓ�_��^[��]� ��D���   �JL�E�P�ыu��P���������D���   ��M�Q�҃�_��^[��]� ���U���SVW3��E��P�M��}��}��E��  �}�}��w��W�M�Q�U�R���T~�����M����7j����t+�u���������D���   ��U�R�Ѓ�_��^[��]� ��D���   �JL�E�P�ыu��P���%�����D���   ��M�Q�҃�_��^[��]� ���U���SVW3��E��P�M��}��}��E��  �}�}���v��W�M�Q�U�R���}�����M����wi��_^��[t��D���   ��U�R�������]Ë�D���   �J<�E�P���]���D���   ��M�Q���E�����]���������������U���SVW3��E��P�M��}��}��E��  �}�}��v��W�M�Q�U�R����|�����M�����h����t��D���   ��U�R�Ѓ�_^3�[��]Ë�D���   �J8�E�P�ы�D�����   ��M�Q�҃�_��^[��]��������������U���SVW3��E��P�M��}��}��E��  �}�}��du��W�M�Q�U�R���4|�����M����h����t-��u��D����   ���^�U�R�Ѓ�_��^[��]� ��D���   �JP�E�P�ы�@�u��D����   �
�F�E�P�у�_��^[��]� �̡�D�PL��  Q��Y��������������U�졨D�PL�E��  ��jPQ�M�Q�ҋ�M�@�A�������]� �������U�졨D�PL�E��  ��j PQ�M�Q�ҋ�M�@�A�������]� �������U���SVW3��E��P�M��}��}��E��  �}�}��t��W�M�Q�U�R����z�����M����f����t-��u��D����   ���^�U�R�Ѓ�_��^[��]� ��D���   �JP�E�P�ы�@�u��D����   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��Ds��W�M�Q�U�R���z�����M�����e����t-��u��D����   ���^�U�R�Ѓ�_��^[��]� ��D���   �JP�E�P�ы�@�u��D����   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��r��W�M�Q�U�R���Ty�����M����7e����t-��u��D����   ���^�U�R�Ѓ�_��^[��]� ��D���   �JP�E�P�ы�@�u��D����   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}���q��W�M�Q�U�R���x�����M����wd����t��D���   ��U�R�Ѓ�_^3�[��]Ë�D���   �J8�E�P�ы�D�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]��E�E�E��P�M��E�   �E��  �q��j�M�Q�U�R����w���M���c����D���   ��U�R�Ѓ�^��]� ���������U����EV��M�E�3�Q�M��E�   �E��  �E�E��p��j�U�R�E�P���w���M��Vc����D���   �
�E�P�у�^��]� ��������U�����D�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��p��j�E�P�M�Q���	w���M���b����D���   ��M�Q�҃�_^��]� ��U�����D�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��o��j�E�P�M�Q���v���M��Qb����D���   ��M�Q�҃�_^��]� ��U�����D�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��o��j�E�P�M�Q���	v���M���a����D���   ��M�Q�҃�_^��]� ��U�����D�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��n��j�E�P�M�Q���u���M��Qa����D���   ��M�Q�҃�_^��]� ��U����EV��M�E�3�Q�M��E�   �E��  �E�E��/n��j�U�R�E�P���u���M���`����D���   �
�E�P�у�^��]� ��������U���SVW3��E��P�M��}��}��E��  �}�}���m��W�M�Q�U�R���t�����M����w`����t-��u��D����   ���^�U�R�Ѓ�_��^[��]� ��D���   �JP�E�P�ы�@�u��D����   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��m��W�M�Q�U�R����s�����M����_����t��D���   ��U�R�Ѓ�_^3�[��]Ë�D���   �J8�E�P�ы�D�����   ��M�Q�҃�_��^[��]��������������U���SVW3��E��P�M��}��}��E��  �}�}��Tl��W�M�Q�U�R���$s�����M����_����t��D���   ��U�R�Ѓ�_^3�[��]Ë�D���   �J8�E�P�ы�D�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U�����D�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��jk��j�E�P�M�Q���Yr���M��!^����D���   ��M�Q�҃�_^��]� ��U����EV��M�E�3�Q�M��E�   �E��  �E�E���j��j�U�R�E�P����q���M��]����D���   �
�E�P�у�^��]� ��������U����EV��M�E�3�Q�M��E�   �E��  �E�E��j��j�U�R�E�P���~q���M��F]����D���   �
�E�P�у�^��]� ��������U�졨D�H���   ]��������������U�졨D�H���   ]�������������̡�D�H���   �⡨D�H���   ��U�졨D�H���   V�u�R�Ѓ��    ^]�����������U�졨D�H���   ]��������������U�졨D�HL�QV�ҋ���u^]á�D�H�U�ER�UP��@  RV�Ѓ���u��D�Q@�BHV�Ѓ�3���^]����������U�졨D�H�U�E��@  R�U�� P�ERP�у�]������U�졨D�H���   ]��������������U�졨D�H�U0�E,R�U(P�E$R�U P�ER�Uj P�ER�UP�ER�UP���   R�Ѓ�0]����������̡�D�PL�BdQ�Ѓ���������������̡�D�PL�BhQ�Ѓ����������������U�졨D�PL�EP�EPQ�Jl�у�]� U�졨D�PL�EPQ��d  �у�]� �U�졨D�PL�EPQ��  �у�]� ̡�D�PL�BtQ�Ѓ����������������U�졨D�PL�EP�EP�EPQ���   �у�]� ���������U�졨D�PL�EP�EP�EPQ�J|�у�]� ������������U���<��DSV��HL�QW�ҋ�3ۉ}�;��w  �M��q����M�E�Qh]  �ȉ]ȉ]Љ]ԉ]؉]��E�   �]��}ĉE�������D���   �PSSW���҅���   ��D�HL�Q W�ҋ���;���   ��    ��D���   �B(���ЍM�Qh�   ���u��ۢ��������   �M�;���   ��D���   ���   S��;�tm��D���   �ȋB<V�Ћ�D���   ���   �E�P�у�;�t��D�B@�HHV�у���;��]����}��M��W���M��������_^[��]� �}���D�B@�HHW�ы�D���   ���   �M�Q�҃��M��jW���M�����_^3�[��]� ������̡�D�PL���   Q�Ѓ������������̡�D�PL���   Q�Ѓ�������������U�졨D�PL�EPQ���   �у�]� ̡�D�PL���   Q�Ѓ�������������U�졨D�PL�EPQ���   �у�]� �U�졨D�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U�E�EVh�� h�� h`� hP� R�Q�UR�UR�UQ�A�$�5�D�vLRP���   Q�Ѓ�,^]� ������������̡�D�PL���   Q�Ѓ�������������U�졨D�PL�EPQ���   �у�]� �U�졨D�PL�EPQ���   �у�]� �U�졨D�PL�EPQ���   �у�]� �U�졨D�PL�EPQ���   �у�]� �U�졨D�PL�EPQ���   �у�]� ̡�D�PL��<  Q�Ѓ�������������U�졨D�PL�EP�EP�EPQ��h  �у�]� ���������U�졨D�PL�EP�EP�EP�EP�EPQ��@  �у�]� �U�졨D�PL�EP�EP�EPQ��D  �у�]� ���������U�졨D�PL�EP�EP�EP�EPQ��H  �у�]� �����U�졨D�HL��$  ]��������������U�졨D�HL��(  ]��������������U�졨D�HL��,  ]�������������̡�D�HL��\  ��U���(��DV3��u؉u܉u��u�u�u�u��E�   �u􋈜   ���   W�ҋ}�E�;�t`;�t\��D�QLjP���   ���ЋM��U�Rh=���M�}��ٝ������D���   ���   �U�R�Ѓ��M؉u��S����_^��]Ë�D���   ���   �E�P�у��M؉u���R��_�   ^��]����������U���(��DV3��u؉u܉u��u�u�u�u��E�   �u􋈜   ���   W�ҋ}�E�;�t`;�t\��D�QLjP���   ���ЋM��U�Rh<���M�}����������D���   ���   �U�R�Ѓ��M؉u��2R����_^��]Ë�D���   ���   �E�P�у��M؉u��R��_�   ^��]���������̋�� h���������h���������̅�t��j�����̡�D�P��l  �ࡨD�P��x  ��U�졨D�P��p  ��V�E�P�ҋuP���
����M��2�����^��]� ��������̡�D�P��t  ��U�졨D�H��d  ]��������������U�졨D�H��  ]�������������̡�D�H��h  ��U�졨D�H��<  ]��������������U�졨D�H���  ]��������������U�졨D�H���  ]��������������U���EV���ht	V��  ����^]� ��������������U��V�u���t��D�QP�B�Ѓ��    ^]���������U�졨D�H��  ]��������������U��E��t�x��u�   ]�3�]������U��E��s�   VW�xW�N  ������u_^]Ã} tWj V�N  ��_������F��D   ^]����������������U���D�E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�M  ������u_^]�Wj V�6N  ��_������F��D   ^]�������������U���D�E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW��L  ������u_^]�Wj V�M  ��_������F��D   ^]�������������U���D�E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�L  ������u_^]�Wj V�6M  ��_������F��D   ^]�������������U���D�E��t#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   VW�xW��K  ������u_^]�Wj V�L  ��_������F��D   ^]���������U���D��tO�} �Et#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËM�UQR�7�����]���U���D�E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�K  ������u_^]�Wj V��K  ��_������F��D   ^]�������������U���D�E��t#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   VW�xW�J  ������u_^]�Wj V�BK  ��_������F��D   ^]���������U���D��tO�} �Et#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËM�UQR�������]���U��M��t.�=�D t�y���A�uP�K  ��]á�D�P�BQ�Ѓ�]�������U��M��t.�=�D t�y���A�uP��J  ��]á�D�P�BQ�Ѓ�]�������U��M��t.�=�D t�y���A�uP�J  ��]á�D�P�BQ�Ѓ�]�������U��M��t.�=�D t�y���A�uP�HJ  ��]á�D�P�BQ�Ѓ�]�������U��M��t.�=�D t�y���A�uP�J  ��]á�D�P�BQ�Ѓ�]�������U��M��t.�=�D t�y���A�uP��I  ��]á�D�P�BQ�Ѓ�]�������U��M��t.�=�D t�y���A�uP�I  ��]á�D�P�BQ�Ѓ�]�������U��M��t.�=�D t�y���A�uP�HI  ��]á�D�P�BQ�Ѓ�]�������U�졨D�H|�]�ࡨD�H|�h   �҃�������������U��V�u���t��D�Q|P�B�Ѓ��    ^]���������U�졨D�P|�EP�EPQ�J�у�]� U�졨D�P|�EP�EPQ�J�у�]� U�졨D�P|�EP�EPQ�J�у�]� U�졨D�P|�EPQ�J�у�]� ����U��Q��D�P�EWP�M�Q�JP�ы�����u_��]� ��D�B��H  SVj �_j S�ы�����u	^[_��]� �M��D�B�U��@TQSVR�Ѓ��> ��^[_��]� ���������������U�졨D�H�Q`VW�}W�ҡ�D�H�U�ADR�Ћ�����t"��D�Q�BpWV�Ћ�D�Q�BV�Ѓ���_^]���������U�졨D�H�Q`V�uV�ҡ�D�H�U�E�I|VRP�у���^]��������������U�졨D�H�Q`VW�}W���E��D�H�U�E��R�UP�ERPQ�I@�$�ы�����t"��D�B�HpWV�ы�D�B�HV�у���_^]���U����13ŉE�V�uW�}�E�0�E�x�   �   ��    ��������
s0�7�D�B��y䡨D�D� �H�Q`W�ҡ�D�H�Adj j��U�RW�ЋM�����_3�^�L=  ��]�������U��� V�uW�}���&  ��   @vp��D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�у��U�Rj0j jj �ǋֱ�JF  �U�E�m�x�]�EQ�E��$P�x�������   ����   ��   v`��D�H�A`�U�R�Ћ�D�Q�Jdj j��E�htP�у��U�Rj0j jj �ǋֱ
��E  �U�E�m�x�]�E�y�����|6��   v,j hp�M��q���mPj0�xj jj �]�E�?���j hl�M��E��P�E�WP�
������uPV�]C����D�Q�Jl�E�P�ы�D�B�Pl�M�Q�҃�_��^��]���������������U��E��u��D�MP�EPQ��E����]��������������̋�3ɉ�H�H�H�U��V��~ W�}u0j j h�Dj�p�������t
W���1����3��F��u_^]� �~ t3�9_��^]� ��D�H<�W�҃�3Ʌ����_�F   ^��]� �����V���F   ��D�H<�Q��3Ʌ����^���������������V��~ t�   ^Ã~ u3�^á�D�H<��AR�ЋN��Q���    �F    ����^����������U����u��D�H�]� ��D�J<�URP�A�Ѓ�]� ���������������U���D��u��D�H�]Ë�D�J<�URP�A�Ѓ�]�U���D��$V��u��D�H�1���D�J<�URP�A�Ѓ�����D�Q�J`�E�SP�ы�D�B�Pp�M�QV�ҡ�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�ы�D�Bj �M�Q�U�R�P$�M�Q�҅���D�H�Al�U�R���Ѓ�4��[t.��D�Q�u�B`V�Ћ�D�Q�Jl�E�P�у���^��]Ë�D�B�M��@,jQ�U�R�Ћ�D�Q�E�M�PQ�J0�E�P�ы�D�B�u�H`V�ы�D�B�Pp�M�VQ�ҡ�D�H�Al�U�R�Ѓ�(��^��]�U���D��$SV��u��D�H�1���D�J<�URP�A�Ѓ�����D�Q�J`�E�P�ы�D�B�Pp�M�QV�ҡ�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�ы�D�Bj �M�Q�U�R�P$�M�Q�҅���D�H�Al�U�R���Ѓ�4��t/��D�Q�u�B`V�Ћ�D�Q�Jl�E�P�у���^[��]Ë�D�B�M��@,jQ�U�R�Ћ�D�Q�E�M�PQ�J0�E�P�ы�D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�Ћ�D�Qj �E�P�M�Q�J$�E�P�ы�D���B�Pl�M�Q���҃�@��t-��D�H�u�Q`V�ҡ�D�H�Al�U�R�Ѓ���^[��]Ë�D�Q�E��R,jP�M�Q�ҡ�D�H�U�E�RP�A0�U�R�Ћ�D�Q�u�B`V�Ћ�D�Q�Jp�E�VP�ы�D�B�Pl�M�Q�҃�(��^[��]�����������U���D��$SV��u��D�H�1���D�J<�URP�A�Ѓ�����D�Q�J`�E�P�ы�D�B�Pp�M�QV�ҡ�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�ы�D�Bj �M�Q�U�R�P$�M�Q�҅���D�H�Al�U�R���Ѓ�4��t/��D�Q�u�B`V�Ћ�D�Q�Jl�E�P�у���^[��]Ë�D�B�M��@,jQ�U�R�Ћ�D�Q�E�M�PQ�J0�E�P�ы�D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�Ћ�D�Qj �E�P�M�Q�J$�E�P�ы�D���B�Pl�M�Q���҃�@��t-��D�H�u�Q`V�ҡ�D�H�Al�U�R�Ѓ���^[��]Ë�D�Q�E��R,jP�M�Q�ҡ�D�H�U�E�RP�A0�U�R�Ћ�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҡ�D�Hj �U�R�E�P�A$�U�R�Ћ�D�Q�Jl���E�P���у�@��t/��D�B�u�H`V�ы�D�B�Pl�M�Q�҃���^[��]á�D�H�U��I,jR�E�P�ы�D�B�M�U�QR�P0�M�Q�ҋu���E�P��������D�Q�Jl�E�P�у���^[��]���������U���D��$SV��u��D�H�1���D�J<�URP�A�Ѓ�����D�Q�J`�E�P�ы�D�B�Pp�M�QV�ҡ�D�H�A`�U�R�Ћ�D�Q�Jdj j��E�h�P�ы�D�Bj �M�Q�U�R�P$�M�Q�҅���D�H�Al�U�R���Ѓ�4��t/��D�Q�u�B`V�Ћ�D�Q�Jl�E�P�у���^[��]Ë�D�B�M��@,jQ�U�R�Ћ�D�Q�E�M�PQ�J0�E�P�ы�D�B�P`�M�Q�ҡ�D�H�Adj j��U�h�R�Ћ�D�Qj �E�P�M�Q�J$�E�P�ы�D���B�Pl�M�Q���҃�@��t-��D�H�u�Q`V�ҡ�D�H�Al�U�R�Ѓ���^[��]Ë�D�Q�E��R,jP�M�Q�ҡ�D�H�U�E�RP�A0�U�R�Ћ�D�Q�J`�E�P�ы�D�B�Pdj j��M�h�Q�ҡ�D�Hj �U�R�E�P�A$�U�R�Ћ�D�Q�Jl���E�P���у�@��t/��D�B�u�H`V�ы�D�B�Pl�M�Q�҃���^[��]á�D�H�U��I,jR�E�P�ы�D�B�M�U�QR�P0�M�Q�҃�j h��M������D�Hj �U�R�E�P�A$�U�R�Ћ�D�Q�Jl���E�P���у����Q�����D�H�U��I,jR�E�P�ы�D�B�M�U�QR�P0�M�Q�ҋu���E�P���e����D�Q�Jl�E�P�у���^[��]���������U�졨D�H<�A]����������������̡�D�H<�Q�����V��~ u>���t��D�Q<P�B�Ѓ��    W�~��t������W�������F    _^��������U���V�E�P��莸����P���#����M��詘����^��]��̃=�D uK��D��t��D�Q<P�B�Ѓ���D    ��D��tV���`���V芗������D    ^������������U���8��D�H�A`S�U�V3�R�]��Ћ�D�Q�JdSj��E�h�P�ы�D�B<�P�M�Q�ҋ�D�H�Al�U�R�Ѓ�;�u^3�[��]�V�M�]��x-  �M�Q�U�R�M���-  ����   W�}�}���   ��D���   �U��ATR�Ћ�����tF��D�Q�J`�E�P���у��U�Rj�E�P��������D�Qj WP�B �Ѓ��E���t�E� ��t��D�Q�Jl�E�P����у���t��D�B�Pl�M�Q����҃��}� u"�E�P�M�Q�M���,  ���7����E�_^[��]ËU��U�_�E�^[��]����������U��E����u��]�VP�M��U,  �EP�M�Q�M��E�    �E    �,  ����   �u�E���tB��t=��u[��D���   �M�PHQ�ҋ�D�Qj VP�B �Ѓ���u-�   ^��]Ë�D���   �E�JTP��VP�V�������uӍUR�E�P�M��,  ���{���3�^��]�V��~ u>���t��D�Q<P�B�Ѓ��    W�~��t��躕��W�������F    _^��������U��E�M�UP��P�EjP�S�����]��������������̸   �����������U��V�u��t���u6�EjP�T�������u3�^]Ë�聄����t���t��U3�;P��I#�^]������̡�D�H\�������U�졨D�H\�AV�u�R�Ѓ��    ^]�������������̡�D�P\�BQ��Yá�D�P\�BQ�Ѓ���������������̡�D�P\�BQ�Ѓ����������������U�졨D�P\�EPQ�J�у�]� ����U�졨D�P\�EP�EPQ�J�у�]� U�졨D�P\�EPQ�J�у�]� ���̡�D�P\�B Q�Ѓ����������������U�졨D�P\�EPQ�J$�у�]� ����U�졨D�P\�EP�EPQ�J(�у�]� U�졨D�P\�EP�EP�EPQ�J,�у�]� ������������U�졨D�P\�EPQ�J4�у�]� ����U�졨D�P\�EPQ�JD�у�]� ����U�졨D�P\�EPQ�JH�у�]� ���̡�D�P\�B8Q�Ѓ����������������U�졨D�P\�EP�EPQ�J<�у�]� U�졨D�P\�EPQ�J@�у�]� ����U���SVW�}��j �ωu��ƨ����D�H\�QV�҃���S��諨��3���~=��I ��D�H\�U�R�U��EP�A,VR�ЋM��Q���x����U�R���m���F;�|�_^[��]� ���������������U���VW�}�E��P��������}� ��   ��D�Q\�B V�Ѓ��M�Q���Ѥ���E���t]S3ۅ�~H�I �UR��赤���E�P��誤���E;E�!����D�Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U��V�u�F��F�����������������]�E��-  �]�����E��������D�Ez��^�P�P�]��������]��E����������N�X�N^�X]�����������U�������P�P��P�P�P�P �P�P�P,�P(�P$�U�M��U��U��U����M��U�P�ɋU��U��U��P�U�H�U��U��M����U��H�M��ɉP�U�U��]��H�M��P�U��]��P$�U��H �M��H(�P,��]�������������U���`�M�A,V�I�A(�I ���I�A(�I�A�I,���I���A�I �A�I���I$���]���E��������Dz�u�؋��������^��]���W���]�A�I,�A�I(�A�I�A�I �A(�I �U��A,�I�]������I$�����I�����e��	���E�������]��A�I�U��A�I�]��A�I,�]��A(�I�U����e��I$�E�������������A�������������]��A�I�A�I �����	�����A�������E��e��I���E�ʍu��ɋ��]��E��e����]��E��e����]����������]��A$�I �A�I,�����]��A,�I�A$�I�����]��A�I�A �I�����]��A(�I�A$�I�����]��A$�I�A(�I�����]��A�I�A�I�   �����]��_^��]�����������U�������P�P��P�P�X���@    �U��U��U��]�M�����M��U��U��P�]�U�P�U��H�M��H�P��]����������U��y t�U��������Au���B�A������Au�B�Y�B�A������Au�B�Y��A������z��Y�B�A������z�B�Y�B�A������z6�B�Y]� �E��Q�P�Q�@�A�Q�A��Q�A�Q�A   ]� ��������U����y ��   ��E�A�]��A�A�]��A�A�]��E��������]�U��E�����]�U�P�M��]��U��P�A� �]��A�`�]�U��A�M��`�E��P�]��M��H��]� ��E�U�V�u��U�U��]�M��P�p�E��P�p^��]� �������������̋�3ɉ�H�H�H�V����t	P��������F�    ��t	P�������F    �F    �F    ^��U��V��W��t	P�������F�    ��t	P�w������}�F    �F    �F    ����   �? ��   �G����   3ɺ   ����j j h�D���Q����������t=� t?�G��t83ɺ   ����j j h�D���Q�������F��u�������_3�^]� �G��F�G��    Q�F�RP�E���F����t�N�W��QPR�xE����_�   ^]� ����������U��SV��3�W;�t	P�j������F�;�t	P�X������^�^�^9]��   �};���   3ɋǺ   ����SSh�D���Q��������;�t>9]tG�]��t@3ɋú   ����j j h�D���Q�������F��u�������_^3�[]� �^�13ɸ   �F�   ����j j h�D���Q�m������F��t���U��    PQR�~�\D���E����t!�N�V��QRP�@D����_^�   []� �F�8_^�   []� 3���A�A�A���U��Q�A�`�
�@�b�	���B�a����]��E���]�������U���|��UV�U��q�<��M��E�    �,  S�]W���  ��Uԋ�UЋM�U̍@�<����}��x�@�E��B�@�����E��}����>��U����]��@�E��������]��@�E��E��E؋E�����E����]ȋEȉE�   ;��  �w����`  �w�����F�B��   �U�P��R�������]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U���P��R���]��E��E��]��E��E��]��E��E��]�����]��B���]��B���]��E����E������E��M������]��E��E������E��ˋU��������]��E��M؉U؋U����ɉU܋U�U����R���]��E��E��]��E��E��]��E��E��]�����]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U��P��R���]��E��E��]��E��E��]��E��E��]���������]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U����]��E��E��]��E��E��]��E��E��]��������U�E��;���   �ۍ�+���@����������]��@���]��@�E����]��E����E������E��M������]��E��E������E����������]��E��M؉E؋E����ɉE܋E�E����]��E��E��]��E��E��]��E��E��]��g�������������������UȋE��UċU��]��M���S�M�Q�U�R�C��������ẺK$�ыP�S(�@�C,������z	�����]��U�E�������z	�����]���U��E�E������E�����   ��������z���]��������z	�����]���U��E�E�������zb�������C(�����C,���]��M��C$���C,�����]ċU��c$�K�S�]ȋEȉC�C�K(�C�K,���]��C�K,�C�K$�   �����������z���]��������z���]��E�E���������   �C,�����C(���]��M��C$�����]ċU��C$���C(�K�ʉS���]ȋEȉC�C(�K�C,�K���]��C,�K�C$�K�M����]ċU��C$�K�C(�K�K�S���]ȋEȉC �{�C(�����C,�������]��M��K$�C,���]ċU��c(�K�S�]ȋEȉC �C�K,�C �K(���]��M��C$�K �C,�K���]ċU��C(�K�C$�K�K�S���]ȋEȉC�M�SQ������U�   �����M������3�3�3���|'�y�����B�U�҉U�U�w����u�U�};�}�Q���U��U�9��E�Ƌu�E����@�����K��@�K���@�K$���]��C��C�@�K���C(�H���]��C��C�@�K ���C,�H�E��E��E����E��]ȋEȉE��E��D��@�����K��@�K���@�K$���]�� �K�C�@�K���C(�H���]�� �K�C�@�K ���C,�H�ẺE����]ԋEЋI���EċE�3��Eȅ���   �F���FU�;���@�E�����K�U���@�K���@�K$���]��C��C�@�K���C(�H���]��C��C�@�K ���@�E��K,���]��E����E������E��U��U��ʉU��E��U����E���E��E��E��E��ʉU��ʉE��������E������]�E�E��]��5����E�_[^��]� �������h�DPh_� �p������������������h�Djh_� �O�������uË@����U��V�u�> t/h�Djh_� �#�������t��U�M�@R�Ѓ��    ^]���U��Vh�Djh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh�Djh_� ����������t�@��t�MQ����^]� 3�^]� �������U��Vh�Djh_� ���i�������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�Djh_� ����������t�@��t�MQ����^]� 3�^]� �������U��Vh�Dj h_� �����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh�Dj$h_� ����������t�@$��t�MQ����^]� 2�^]� �������Vh�Dj(h_� ���\�������t�@(��t��^��3�^������Vh�Dj,h_� ���,�������t�@,��t��^��3�^������U��Vh�Dj0h_� �����������t�@0��t�MQ����^]� 3�^]� �������U��Vh�Dj4h_� ����������t�@4��t�M�UQR����^]� ���^]� ��Vh�Dj8h_� ���|�������t�@8��t��^��3�^������U��Vh�Dj<h_� ���I�������t�@<��t�MQ����^]� ��������������U��Vh�Dj@h_� ���	�������t�@@��t�MQ����^]� ��������������U��Vh�DjDh_� �����������t�@D��t�MQ����^]� 3�^]� �������U��Vh�DjHh_� ����������t�@H��t�MQ����^]� ��������������Vh�DjLh_� ���L�������t�@L��t��^��3�^������Vh�DjPh_� ����������t�@P��t��^��^��������Vh�DjTh_� �����������t�@T��t��^��^��������Vh�DjXh_� ����������t�@X��t��^��^��������U��Vh�Dj\h_� ����������t�@\��t�M�UQR����^]� 3�^]� ���U��Vh�Dj`h_� ���I�������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�Djdh_� ���	�������t�@d��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh�Djhh_� ����������t�@h��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�Djlh_� ���i�������t�@l��t�M�UQR����^]� 3�^]� ���U��Vh�Djph_� ���)�������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh�Djth_� �����������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�Djxh_� ����������t�@x��t�MQ����^]� 3�^]� �������U��Vh�Dj|h_� ���i�������t�@|��t�M�UQR����^]� 3�^]� ���U��Vh�Dh�   h_� ���&�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�Dh�   h_� �����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U���X��A�U�V�U��]����z  S��E��EW����������O  ���������U�r�z�
�R;��4v���I�$��4����R����   �]��F�a�]��F�a�]���!�]��B�a�]��B�a�]��E����E������E����E����������]��E������E������������]��������]��E��E��]��E��E��]��E��   �]��F�a�]��F�a����]���!�]��B�a�]��B�a�]��E����E������E����E����������]��E������E������������]��������]��E��E��]��E��E��]��E��E��]����m������_[�u�E�PV���������^��]� U���$V��M�������F����   �6S�]W�u��E���$    ���������t[��%�����E�M܋���@��P�����F�@��R�M�������~���Q�M�������v;�t�v��P�M�������u����m��u�u�_[�M�UQR�M��v���^��]� ��������������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$�x+�E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��+(+;+O+c+����U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V����t	P�1������F�    ��t	P�������F    �F    �F    ^��U��3�V���F�F�F�EP�D�����^]� �������������U��EVP���!�����^]� ����������U��SV��W3�;�t	P�������F�>;�t	P�������]�~�~�~;�to3ɋú   ����WWh�D���Q�&��������tG�}��tI3ɋǺ   ����j j h�D���Q��������F��u���t	P�������    _^3�[]� �~_�^^�   []� �����������U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��3�V��W�}��F�F�F�Gj;Gu2j������tY�����O�H�G��B�N_���   ^]� j�f�����t'�����W�Q��O�H��G�B�N�   _��^]� ���U��E��u�E�M��D��D�   ]� �����������U��EHV����   �$��/�   ^]á�D@��D��uQ�EP������=�*  }�����^]Ëu��t�j j h�Dj�j������t ����j����D��tV���_m���   ^]���D    �   ^]ËM�UQR�(���������H^]�^]�C
���-�Du.��
��������D��t���k��V�9j������D    �   ^]Ã��^]Ë��.f/m/�.�/K/����U�졨D���   �BXQ�Ѓ���u]� ��D���   �M�RQ�MQP�҃�]� U�졨D���   �BXQ�Ѓ���u]� ��D���   �M�R8Q�MQP�҃�]� U��EV��j ���D�Qj j P���   �ЉF����^]� ��DVj ��H����   j j R�Ѓ��F^�������������U��V��F��u^]� ��D�Q�MP�EP�Q���   P�у��F�   ^]� �9H�X1�\1 ?�`1�>�d1?�h1v>�l1�p1�G�t1�>�x1�=�|1�=Ë�U�������  �} ��Dt�  ��]�;1u���  ��U��EVW��u|P��)  Y��u3��  ��  ��u��)  ���g)  � �a� (  ��D�A"  ��}�e  ���K'  ��| ��$  ��|j ��  Y��u��D�   �\$  ��3�;�u19=�D~���D9=lHu�!  9}u{�/$  �  �Y)  �j��uY�  h  j�  ��YY;��6���V�5�1�54H�  Y�Ѕ�tWV��  YY� �N���V�  Y�������uW�y  Y3�@_^]� jh�!��*  ����]3�@�E��u9�D��   �e� ;�t��u.����tWVS�ЉE�}� ��   WVS�r����E����   WVS�^����E��u$��u WPS�J���Wj S�B�������tWj S�Ѕ�t��u&WVS�"�����u!E�}� t����tWVS�ЉE��E������E���E��	PQ��)  YYËe��E�����3��**  Ë�U��}u��+  �u�M�U�����Y]� �U��WV�u�M�}�����;�v;���  ��   r�=�_ tWV����;�^_u^_]�,  ��   u������r*��$�D5��Ǻ   ��r����$�X4�$�T5��$��4�h4�4�4#ъ��F�G�F���G������r���$�D5�I #ъ��F���G������r���$�D5�#ъ���������r���$�D5�I ;5(5 5555 5�4�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�D5��T5\5h5|5�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��6�����$��6�I �Ǻ   ��r��+��$��5�$��6��56@6�F#шG��������r�����$��6�I �F#шG�F���G������r�����$��6��F#шG�F�G�F���G�������V�������$��6�I �6�6�6�6�6�6�6�6�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��6���6�677�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̃=�_ t-U�������$�,$�Ã=�_ t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�Ë�Q���B*  YË�U��V��������EtV����Y��^]� ��U��� S3�9]u�R=  SSSSS�    ��<  ������N�E;�t�V�u�E��u�E��u�E�P�E�����E�B   ��/  ���M��x�E����E�PS�-  YY��^[�Ë�U���uj �u�u�m�����]�jh�!��$  �e� �u;5�_w"j�r>  Y�e� V�yF  Y�E��E������	   �E���$  �j�m=  YË�U��V�u�����   SW�= �=�I u��,  j�+  h�   �G  YY��_��u��t���3�@P���uV�S���Y��u��uF�����Vj �5�I�׋؅�u.j^9Nt�u�H  Y��t�u�{�����;  �0��;  �0_��[�V�H  Y��;  �    3�^]���̋T$�L$��ti3��D$��u��   r�=�_ t��H  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh�!�:#  �u��tu�=�_uCj��<  Y�e� V�=  Y�E��t	VP�$=  YY�E������   �}� u7�u�
j��;  Y�Vj �5�I� ��u��:  ��� P�r:  �Y��"  ��������̀�@s�� s����Ë������������Ë�U��QSVW�5a�{  �5a���}��k  ��YY;���   ��+ߍC��rwW�H  ���CY;�sH�   ;�s���;�rP�u��J  YY��u�G;�r@P�u��4  YY��t1��P�4��  Y�a�u�x  ���V�m  Y�a�EY�3�_^[�Ë�Vjj �  ��V�F  ���a�a��ujX^Ã& 3�^�jh"�!  �  �e� �u�����Y�E��E������	   �E��!  ��}  Ë�U���u���������YH]�̃��$�mJ  �   ��ÍT$�J  R��<$�D$tQf�<$t��I  �   �u���=�D �CJ  �   �P1�@J  �  �u,��� u%�|$ u���I  �"��� u�|$ u�%   �t����-P5�   �=�D ��I  �   �P1��H  ZË�U��EV���F ��uc��  �F�Hl��Hh�N�;�;t��:�Hpu�ET  ��F;�9t�F��:�Hpu�L  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P��U  ��e�F�P�T  ��Yu��P��U  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�U  �M��E��M��H��EP�U  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�Y  @PV�V�V  ��^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M�������3�;�u+�-6  j_VVVVV�8�5  ���}� t�E��`p����!  9uv�9u~�E�3���	9Ew	��5  j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h�SV��X  ��3ۅ�tSSSSS��3  ���N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�TNt�90uj�APQ�T  ���}� t�E��`p�3�_^[�Ë�U���,�13ŉE��ESVW�}j^V�M�Q�M�Q�p�0�Z  3ۃ�;�u�4  SSSSS�0�.4  �����o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q�4X  ��;�t���u�E�SP�u��V�u��������M�_^3�[�����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �C���9}}�}�u;�u+�3  j^WWWWW�0�A3  ���}� t�E�`p����  9}vЋE��� 9Ew	�z3  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�%E  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� ��X  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �X  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V������u�E�8 u���} �4����$�p���WF�X  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP��V  0�F�U�����;�u��|��drj jdRP��V  0��U�F����;�u��|��
rj j
RP�V  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N�������u-�W0  j^�03�PPPPP��/  ���}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V��������}� t�E��`p�3�_^[�Ë�U���,�13ŉE��ESVW�}j^V�M�Q�M�Q�p�0��T  3ۃ�;�u�H/  SSSSS�0��.  �����Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P��R  ��;�t���u�E�SV�u���`������M�_^3�[�����Ë�U���0�13ŉE��ESV�uWj_W�M�Q�M�Q�p�0�T  3ۃ�;�u�.  SSSSS�8�.  �����   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW�4R  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[������Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3���X1�6�  ��Y���(r�_^Ë�Vh   h   3�V��S  ����tVVVVV�P+  ��^Ë�U������]����]��E��u��M��m��]����]�����z3�@��3���h�� ��th�P� ��tj ���������U���(  �F�F�F�F�5 F�=�Ef�(Ff�Ff��Ef��Ef�%�Ef�-�E�� F�E �F�E�F�E�$F�������`E  �F�E�E	 ��E   �1������� 1�������0 �XEj�S  Yj �, h�( �=XE uj��R  Yh	 ��$ P�  �Ë�U��V�5�1�58 �օ�t!��1���tP�5�1���Ѕ�t���  �'� V�4 ��uV�  Y��thP� ��t�u�ЉE�E^]�j ����YË�U��V�5�1�58 �օ�t!��1���tP�5�1���Ѕ�t���  �'� V�4 ��uV�   Y��th<P� ��t�u�ЉE�E^]��< � ��V�5�1�8 ����u�50H�e���Y��V�5�1�@ ��^á�1���tP�58H�;���Y�Ѓ�1���1���tP�D ��1��*  jh0"�  � V�4 ��uV�a  Y�E�u�F\�3�G�~��t$hP� �Ӊ��  h<�u��Ӊ��  �~pƆ�   CƆK  C�Fh�5j�O+  Y�e� �vh�H �E������>   j�.+  Y�}��E�Fl��u��;�Fl�vl��C  Y�E������   �  �3�G�uj�*  Y�j�*  YË�VW� �5�1�������Ћ���uNh  j��  ��YY��t:V�5�1�54H�����Y�Ѕ�tj V�����YY� �N���	V�}���Y3�W�L _��^Ë�V��������uj�>  Y��^�jhX"�  �u����   �F$��tP�0���Y�F,��tP�"���Y�F4��tP����Y�F<��tP����Y�F@��tP�����Y�FD��tP�����Y�FH��tP�����Y�F\=�tP�����Yj��)  Y�e� �~h��tW�P ��u���5tW����Y�E������W   j�)  Y�E�   �~l��t#W��B  Y;=�;t���:t�? uW��@  Y�E������   V�F���Y��  � �uj�W(  YËuj�K(  YË�U��=�1�tK�} u'V�5�1�58 �օ�t�5�1�5�1���ЉE^j �5�1�54H����Y���u�x�����1���t	j P�@ ]Ë�VW� V�4 ��uV�R  Y�����^  �5 hlW��h`W�,H��hTW�0H��hLW�4H�փ=,H �5@ �8Ht�=0H t�=4H t��u$�8 �0H�D �,HK�54H�8H�< ��1�����   �50HP�օ���   �_  �5,H�����50H�,H�����54H�0H�����58H�4H�u������8H�&  ��teh�L�5,H�����Y�У�1���tHh  j�   ��YY��t4V�5�1�54H����Y�Ѕ�tj V�y���YY� �N��3�@��$���3�_^Ë�U��VW3��u�������Y��u'9<HvV�T ���  ;<Hv��������uʋ�_^]Ë�U��VW3�j �u�u�L  ������u'9<HvV�T ���  ;<Hv��������uË�_^]Ë�U��VW3��u�u�UM  ��YY��u,9Et'9<HvV�T ���  ;<Hv��������u���_^]Ë�U��W��  W�T �u�4 ���  ��`�  w��t�_]Ë�U����  �u�  �5�1�D���h�   �Ѓ�]Ë�U��h��4 ��thxP� ��t�u��]Ë�U���u�����Y�u�X �j�%  Y�j��$  YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=� th���N  Y��t
�u��Y�B���h@h,����YY��uBhD[������ �$(�c����=a Ytha�rN  Y��tj jj �a3�]�jh�"�  j��$  Y�e� 3�C9pH��   �lH�E�hH�} ��   �5a�����Y���}؅�tx�5a����Y���u܉}�u����u�;�rW����9t�;�rJ�6��������������5a�~������5a�q�����9}�u9E�t�}�}؉E����u܋}��hP�D�_���YhX�T�O���Y�E������   �} u(�pHj��"  Y�u�����3�C�} tj��"  Y��7
  Ë�U��j j�u�������]�jj j ������Ë�V������V�k.  V�P  V�   V�M  V��O  V��M  V�  V��M  h�S������$��1^�jTh�"�r	  3��}��E�P�h �E�����j@j ^V�&���YY;��  � `�5�_��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@� `��   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M��� `���_ ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=�_|���=�_�e� ��~m�E����tV���tQ��tK�uQ�d ��t<�u���������4� `�E� ���Fh�  �FP�}N  YY����   �F�E�C�E�9}�|�3ۋ���5 `����t���t�N��r�F���uj�X�
��H������P�` �����tC��t?W�d ��t4�>%�   ��u�N@�	��u�Nh�  �FP��M  YY��t7�F�
�N@�����C���g����5�_�\ 3��3�@Ëe��E���������p  Ë�VW� `�>��t1��   �� t
�GP�l ���@   ;�r��6�����& Y���� a|�_^Ã=a u��7  V�5�DW3���u����   <=tGV�A  Y�t���u�jGW�n�����YY�=PH��tˋ5�DS�BV�lA  ��C�>=Yt1jS�@���YY���tNVSP��A  ����t3�PPPPP�  �����> u��5�D������%�D �' � a   3�Y[_^��5PH������%PH ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF��L  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#��K  Y��t��M�E�F��M��E����K  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9au�l5  h  �xHVS�|I�p �a�5`H;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�q�����Y;�t)�U��E�P�WV�}�������E���H�DH�5HH3�����_^[�Ë�U�졀I��SV�5� W3�3�;�u.�֋�;�t��I   �#� ��xu
jX��I���I����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5� SSS+�S��@PWSS�E��։E�;�t/P����Y�E�;�t!SS�u�P�u�WSS�օ�u�u�����Y�]��]�W�| ���\��t;�u��x ��;��r���8t
@8u�@8u�+�@P�E��0�����Y;�uV�t �E����u�VW�������V�t ��_^[�Ë�V��!��!W��;�s���t�Ѓ�;�r�_^Ë�V��!��!W��;�s���t�Ѓ�;�r�_^Ë�U��3�9Ej ��h   P�� ��I��u]�3�@��_]Ã=�_uWS3�9�_W�= ~3V�5�_��h �  j �v��� �6j �5�I�׃�C;�_|�^�5�_j �5�I��_[�5�I�� �%�I �Ë�U��QQV�G��������F  �V\��1W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ��1�=�1���;�}$k��~\�d9 �=�1��1B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]��h�]d�5    �D$�l$�l$+�SVW�11E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s351W��E� �E�   �{���t�N�38�I����N�F�38�9����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���HG  �E���|@G�E��؃��u΀}� t$����t�N�38������N�V�3:�����E�_^[��]��E�    �ɋM�9csm�u)�=�_ t h�_��A  ����t�UjR��_���M��F  �E9Xth1W�Ӌ���F  �E�M��H����t�N�38�3����N�V�3:�#����E��H���F  �����9S�R���h1W���F  ������U����1�e� �e� SW�N�@��  ��;�t��t	�У 1�`V�E�P�� �u�3u��� 3�� 3��� 3��E�P�� �E�3E�3�;�u�O�@����u������51�։5 1^_[��U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]�jh�"�����e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E��
���Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[��������_3��jh�"�I���j��  Y�e� �u�N��t/��I��I�E��t9u,�H�JP�����Y�v�����Y�f �E������
   �8���Ë���j��  Y�����̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�U���(  �13ŉE���1Vtj
��   Y��>  ��tj��>  Y��1��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P���������������(�����0���j ǅ����  @��������,����, ��(���P�( j�Q���̋�U��QQS�]VW3�3��}�;��1t	G�}���r���w  j�4D  Y���4  j�#D  Y��u�= E�  ���   �A  h��  S��IW�A4  ����tVVVVV�  ��h  ��IVj ��J �p ��u&h�h�  V��3  ����t3�PPPPP��  ��V�X3  @Y��<v8V�K3  ��;�j��Lh�+�QP�B  ����t3�VVVVV�  ���3�h�SW�B  ����tVVVVV�m  ���E��4��1SW��A  ����tVVVVV�H  ��h  hxW�i@  ���2j��` ��;�t$���tj �E�P�4��1�6�2  YP�6S�� _^[��j�B  Y��tj�B  Y��u�= Euh�   �)���h�   ����YYË�U��E��L]Ë�U��QV�uV��N  �E�FY��u�!  � 	   �N ����/  �@t�  � "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�L  �� ;�t�L  ��@;�u�u�?L  Y��uV��K  Y�F  W��   �F�>�H��N+�I;��N~WP�u��J  ���E��M�� �F����y�M���t���t����������� `���1�@ tjSSQ�HB  #����t%�F�M��3�GW�EP�u�pJ  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u�O  �8*u�ϰ?�d����} �^[]Ë�U���x  �13ŉE�S�]V�u3�W�}�u�������������������������������������������������������������G�����u5��  �    3�PPPPP�M  �������� t
�������`p������
  �F@u^V�;L  Y��1���t���t�ȃ�������� `����A$u����t���t�ȃ������ `����@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw�������3��3�3�����j��Y������;���	  �$��s��������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�������K  Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u��2������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P�bI  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ��2������P�i*  Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7����������F  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V�����������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5p1�����Y�Ћ���������   t 9�����u������PS�5|1�����Y��YY������gu;�u������PS�5x1����Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW��E  ��0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u��2�������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF��C  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t����������������� Y���������������t������������������������� t
�������`p��������M�_^3�[豽���Ð�k�i j^j�j�j�j)l��U��E��L]Ë�U���(  �13ŉE������� SjL������j P������������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������0 j ���, ��(���P�( ��u��uj��'  Yh ��$ P�  �M�3�[�Y����Ë�U���5�L�e���Y��t]��j�'  Y]������U��E3�;͸2tA��-r�H��wjX]Ëͼ2]�D���jY;��#���]��������u� 4Ã���������u�$4Ã�Ë�U��V������MQ�����Y�������0^]Ë�VW3���L�<�,4u��(4�8h�  �0���.  YY��tF��$|�3�@_^Ã$�(4 3����S�l V�(4W�>��t�~tW��W�����& Y����H5|ܾ(4_���t	�~uP�Ӄ���H5|�^[Ë�U��E�4�(4�� ]�jh #�����3�G�}�3�9�Iu�T���j����h�   �����YY�u�4�(49t���nj�N���Y��;�u�����    3��Qj
�Y   Y�]�9u,h�  W�-  YY��uW�<���Y�o����    �]���>�W�!���Y�E������	   �E������j
�(���YË�U��EV�4�(4�> uP�"���Y��uj�����Y�6�� ^]Ë�U���_��_k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �N����   ��_�5� h @  ��H� �  SQ�֋�_�N�   ���	P�N�@��_����    �N�@�HC�N�H�yC u	�`��N�x�ueSj �p�֡N�pj �5�I� ��_�Nk���_+ȍL�Q�HQP�  �E����_;Nv�m��_��_�E�N�=�_[_^�á�_V�5�_W3�;�u4��k�P�5�_W�5�I�� ;�u3��x��_�5�_��_k�5�_h�A  j�5�I� �F;�t�jh    h   W�� �F;�u�vW�5�I� 뛃N��>�~��_�F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�� ��u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U�����_�Mk��_������M���SI�� VW}�����M���������3���U���_����S�;#U�#��u
���];�r�;�u��_��S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1��_�	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t��_�C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;Nu�M�;�_u�%N �M���B_^[�Ë�U��E�N]Ë�U���5N�2���Y��t�u��Y��t3�@]�3�]�U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh #�(���3��]3�;���;�u�����    WWWWW����������S�=�_u8j����Y�}�S�����Y�E�;�t�s���	�u���u��E������%   9}�uSW�5�I�� ����������3��]�u�j�q���Y�̀zuf��\���������?�f�?f��^���٭^����l5�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����l5�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����d5���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-P5��p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�/4  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��`�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��������������|�����   s�����������������t�����   v��������U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP蝱��3��ȋ��~�~�~����~�����5���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �13ŉE�SW������P�v�� �   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R�ڰ����C�C��u�j �v�������vPW������Pjj �8  3�S�v������WPW������PW�vS��5  ��DS�v������WPW������Ph   �vS�5  ��$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[�a�����jh@#�q�����������:�Gpt�l t�wh��uj �����Y�������j�����Y�e� �wh�u�;5�9t6��tV�P ��u���5tV�Ư��Y��9�Gh�5�9�u�V�H �E������   뎋u�j����YË�U���S3�S�M��/����N���u�N   �� 8]�tE�M��ap��<���u�N   �� �ۃ��u�E��@�N   ��8]�t�E��`p���[�Ë�U��� �13ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9��9��   �E��0=�   r����  �p  ����  �d  ��P�� ���R  �E�PW�� ���3  h  �CVP�����3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP賭���M��k�0�u����9�u��*�F��t(�>����E����9D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C���9Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95N�X�������M�_^3�[�\�����jh`#�l����M��诿�����}�������_h�u�u����E;C�W  h   �����Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�P ��u�Fh=�5tP袬��Y�^hS�=H ���Fp��   ��:��   j�u���Y�e� �C�$N�C�(N�C�,N3��E��}f�LCf�EN@��3��E�=  }�L���7@��3��E�=   }��  ���8@���5�9�P ��u��9=�5tP����Y��9S���E������   �0j�����Y��%���u ���5tS賫��Y������    ��e� �E��$���Ã=a uj��V���Y�a   3�Ë�U��SV�u���   3�W;�to=�>th���   ;�t^9uZ���   ;�t9uP�:������   �#4  YY���   ;�t9uP�������   �3  YY���   �������   �����YY���   ;�tD9u@���   -�   P�ժ�����   ��   +�P�ª�����   +�P贪�����   詪�������   �=(>t9��   uP�1  �7肪��YY�~P�E   ���:t�;�t9uP�]���Y9_�t�G;�t9uP�F���Y���Mu�V�7���Y_^[]Ë�U��SV�5H W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��:t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5P W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��:t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Å�t7��t3V�0;�t(W�8�����Y��tV�E����> Yu���:tV�Y���Y��^�3��jh�#�����L�����:�Fpt"�~l t�5����pl��uj �z���Y�������j����Y�e� �Fl�=�;�i����E��E������   ��j�~���Y�u�Ë�U����u�M������E����   ~�E�Pj�u�>2  ������   �M�H���}� t�M��ap��Ë�U��=0N u�E�x;�A��]�j �u����YY]Ë�U���SV�u�M��q����]�   ;�sT�M胹�   ~�E�PjS�1  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P��#  YY��t�Ej�E��]��E� Y��X���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P��+  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=0N u�E�H���w�� ]�j �u�����YY]Ë�U���(�13ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P�;  �E�E�VP�1  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�����Ë�U���(�13ŉE�SV�uW�u�}�M��w����E�P3�SSSSW�E�P�E�P�;  �E�E�VP�5  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�o����������������U��WV�u�M�}�����;�v;���  ��   r�=�_ tWV����;�^_u^_]�B�����   u������r*��$�����Ǻ   ��r����$����$�����$�����ԕ��#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I {�h�`�X�P�H�@�8��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$� ������$�З�I �Ǻ   ��r��+��$�$��$� ��4�X����F#шG��������r�����$� ��I �F#шG�F���G������r�����$� ���F#шG�F�G�F���G�������V�������$� ��I ԗܗ���������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$� ���0�8�H�\��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��MS3�VW;�t�};�w�[���j^�0SSSSS����������0�u;�u��ڋъ�BF:�tOu�;�u�� ���j"Y�����3�_^[]Ë�U��MSV�u3�W�y;�u�����j^�0SSSSS�}��������   9]v݋U;ӈ~���3�@9Ew����j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�a���@PWV�������3�_^[]Ë�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���H���u��P������Ɂ���  �P���t�M�_^f�H[�Ë�U���0�13ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��c;  �uЉC�E։�EԉC�E�P�uV������$��t3�PPPPP�������M�_�s^��3�[��������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j詴��YË�U��E�M%����#�V������t1W�}3�;�tVV�6D  YY������j_VVVVV�8�O�������_��uP�u��t	�D  ����C  YY3�^]Ã%�_ �jh�#�����M3�;�v.j�X3���;E�@u�^����    WWWWW�������3���   �M��u;�u3�F3ۉ]���wi�=�_uK������u�E;�_w7j�����Y�}��u�����Y�E��E������_   �]�;�t�uWS�&�����;�uaVj�5�I� ��;�uL9=Nt3V�z���Y���r����E;��P����    �E���3��uj�o���Y�;�u�E;�t�    ��輿���jh�#�j����]��u�u�Κ��Y��  �u��uS����Y�  �=�_��  3��}�����  j�����Y�}�S����Y�E�;���   ;5�_wIVSP���������t�]��5V����Y�E�;�t'�C�H;�r��PS�u�����S�����E�SP�������9}�uH;�u3�F�u������uVW�5�I� �E�;�t �C�H;�r��PS�u�踔��S�u��������E������.   �}� u1��uF������uVSj �5�I�� ����u�]j�	���YË}����   9=Nt,V�����Y������������9}�ul��� P����Y��_����   �����9}�th�    �q��uFVSj �5�I�� ����uV9Nt4V�e���Y��t���v�V�U���Y�����    3��ɽ����q����|�����u�c������ P�����Y��������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�#h�]d�    P��SVW�11E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh $������>����@x��t�e� ���3�@Ëe��E������x��������h���E���Y�XNË�U��E�\N�`N�dN�hN]Ë�U��E��1V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5dN�Y���Y�j h $�K���3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�������}؅�u����a  �\N�\N�`�w\���]���������Z�Ã�t<��t+Ht������    3�PPPPP�T�����뮾dN�dN��`N�`N�
�hN�hN�E�   P蕧���E�Y3��}���   9E�uj舰��9E�tP�&���Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.��1�M܋�1��1�9M�}�M�k��W\�D�E����������E������   ��u�wdS�U�Y��]�}؃}� tj ����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3�����Ë�U��E�pN]Ë�U��E�tN]�jh@$�}����e� �u�u�� �E��/�E� � �E�3�=  �����Ëe�}�  �uj�L �e� �E������E��o���Ë�U����u�M�耘���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]���SVW�T$�D$�L$URPQQhd�d�5    �13ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C��?  �   �C��?  �d�    ��_^[ËL$�A   �   t3�D$�H3�����U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�'?  3�3�3�3�3���U��SVWj j h�Q�U  _^[]�U�l$RQ�t$������]� ��U���SVW�P����e� �=�N ����   h��� �����*  �5 h�W�օ��  P蚣���$�W��N��P腣���$|W��N��P�p����$`W��N��P�[���Y��N��thHW��P�C���Y��N��N;�tO9�NtGP衣���5�N��蔣��YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9��N;�t0P�Q���Y��t%�ЉE���t��N;�tP�4���Y��t�u��ЉE��5�N����Y��t�u�u�u�u����3�_^[�Ë�U��ES3�VW;�t�};�w�����j^�0SSSSS�_��������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u�����j"Y����3�_^[]Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w�M���j^�0SSSSS�����������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x���������j"Y���낋�U��MV3�;�|��~��u��D�(��D��D�����VVVVV�    � ��������^]Ë�U��E��t���8��  uP�)���Y]Ë�U��QQ�EV�u�E��EWV�E�� =  ���Y;�u�4���� 	   �ǋ��J�u�M�Q�u�P�� �E�;�u� ��t	P�&���Y�ϋ����� `�����D0� ��E��U�_^��jh`$�۳������u܉u��E���u������  ����� 	   �Ƌ���   3�;�|;�_r!�����8����� 	   WWWWW�������ȋ����� `��������L1��u&�`����8�F���� 	   WWWWW�������������[P�\<  Y�}���D0t�u�u�u�u�������E܉U�������� 	   � ����8�M���M���E������   �E܋U�������u�<  YË�U���  �>  �13ŉE��EV3���4�����8�����0���9uu3���  ;�u'�����0�t���VVVVV�    �����������  SW�}�����4� `�����ǊX$�����(�����'�����t��u0�M����u&�%���3��0�	���VVVVV�    �������C  �@ tjj j �u�~������u�i  Y����  ��D���  �����@l3�9H�������P��4�� ����� ���`  3�9� ���t���P  �� ��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P�
  Y��t:��4���+�M3�@;���  j��@���SP�<  �������  C��D����jS��@���P�<  �������  3�PPj�M�Qj��@���QP�����C��D����� �����\  j ��<���PV�E�P��(���� �4�� ���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4�� ����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@����9  Yf;�@����h  ��8����� ��� t)jXP��@����p9  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4�� ���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4�� ���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �� ��;���   j ��,���P��+�P��5����P��(���� �4�� ��t�,���;���� ��@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0�� ��t��,�����@��� ��8����� ��@�����8��� ul��@��� t-j^9�@���u������ 	   �����0�?��@�������Y�1��(�����D@t��4����8u3��$�����    ������  ������8���+�0���_[�M�3�^�����jh�$菫���E���u�����  �m���� 	   ����   3�;�|;�_r!�_����8�E���� 	   WWWWW��������ɋ����� `��������L1��t�P�@4  Y�}���D0t�u�u�u�.������E�������� 	   ������8�M���E������	   �E�������u�4  YË�U����Nh   �:���Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u�W���� 	   3�]�V3�;�|;�_r�9���VVVVV� 	   �������3���ȃ����� `���D��@^]ø�;á�_Vj^��u�   �;�}�ƣ�_jP躜��YY��O��ujV�5�_衜��YY��O��ujX^�3ҹ�;���O��� ���� >|�j�^3ҹ�;W������ `����������t;�t��u�1�� B��<|�_3�^��7  �=hH t�c5  �5�O�����YË�U��V�u��;;�r"�� >w��+�����Q������N �  Y�
�� V�� ^]Ë�U��E��}��P�����E�H �  Y]ËE�� P�� ]Ë�U��E��;;�r= >w�`���+�����P�y���Y]Ã� P�� ]Ë�U��M���E}�`�����Q�J���Y]Ã� P�� ]Ë�U��EV3�;�u�<���VVVVV�    �Ŀ���������@^]á1��3�9�N����Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�ƿ��j^SSSSS�0�O��������V�u�M������E�9X��   f�E��   f;�v6;�t;�vWSV�ȃ�����s���� *   �h���� 8]�t�M��ap�_^[��;�t2;�w,�H���j"^SSSSS�0�Ѿ����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�� ;�t9]�^����M;�t���� ��z�D���;��g���;��_���WSV�������O�����U��j �u�u�u�u�|�����]Ë�U����u�M������E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]��V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U���VW�u�M�� ����E�u3�;�t�0;�u,�r���WWWWW�    ��������}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP��  �M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&�ѻ���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u90Nuh�;�P������]Ë�S��QQ�����U�k�l$���   �13ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|�����3  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�3  ��h��  ��x�����5  �>YYt�=h@ uV�5  Y��u�6�T5  Y�M�_3�^��u����]��[Ë�U����13ŉE�SV3�W��9�Nu8SS3�GWhh   S�� ��t�=�N�� ��xu
��N   9]~"�M�EI8t@;�u�����E+�H;E}@�E��N����  ;���  ����  �]�9] u��@�E �5� 3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�)  ��;�t� ��  �P�w|��Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5� SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�Y(  ��;�tj���  ���P�{��Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�� ��t"SS9]uSS��u�u�u�VS�u �� �E�V�^���Y�u��U����E�Y�Y  �]�]�9]u��@�E9] u��@�E �u�"4  Y�E���u3��!  ;E ��   SS�MQ�uP�u �@4  ���E�;�tԋ5� SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�C'  ��;�t����  ���P�z��Y;�t	� ��  �����3�;�t��u�SW�J{�����u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��3  ���u������#u�W�3���Y��u�u�u�u�u�u�� ��9]�t	�u��O{��Y�E�;�t9EtP�<{��Y�ƍe�_^[�M�3��Qr���Ë�U����u�M���}���u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap��Ë�U��QQ�13ŉE���NSV3�W��;�u:�E�P3�FVhV�� ��t�5�N�4� ��xu
jX��N���N����   ;���   ����   �]�9]u��@�E�5� 3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�\%  ��;�t� ��  �P�x��Y;�t	� ��  ���؅�ti�?Pj S�hy����WS�u�uj�u�օ�t�uPS�u�� �E�S�o����E�Y�u3�9]u��@�E9]u��@�E�u�C1  Y���u3��G;EtSS�MQ�uP�u�k1  ����;�t܉u�u�u�u�u�u�� ��;�tV�=y��Y�Ǎe�_^[�M�3��Rp���Ë�U����u�M���{���u$�M��u �u�u�u�u�u�������}� t�M��ap��Ë�U��V�u����  �v��x���v��x���v�x���v�x���v�x���v�x���6�x���v �x���v$�x���v(�x���v,�~x���v0�vx���v4�nx���v�fx���v8�^x���v<�Vx����@�v@�Kx���vD�Cx���vH�;x���vL�3x���vP�+x���vT�#x���vX�x���v\�x���v`�x���vd�x���vh��w���vl��w���vp��w���vt��w���vx��w���v|��w����@���   ��w�����   �w�����   �w�����   �w�����   �w�����   �w�����   �w�����   �xw�����   �mw�����   �bw�����   �Ww����,^]Ë�U��V�u��t5�;�>tP�4w��Y�F;�>tP�"w��Y�v;5�>tV�w��Y^]Ë�U��V�u��t~�F;�>tP��v��Y�F;�>tP��v��Y�F;�>tP��v��Y�F; ?tP�v��Y�F;?tP�v��Y�F ;?tP�v��Y�v$;5?tV�v��Y^]�����U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U���S�u�M��x���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�[���YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�8����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���58?N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�4?��+8?;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�58?N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��<?A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;0?�<?��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�0?�D?�3�@�   �D?�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+<?��M���Ɂ�   �ً@?]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5P?N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�L?��+P?;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5P?N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��T?A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;H?�T?��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�H?�\?�3�@�   �\?�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+T?��M���Ɂ�   �ًX?]���@u�M�U�Y��
�� u�M�_[�Ë�U���|�13ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u蓥��SSSSS�    ������3��N  �U�U��< t<	t<
t<uB��0�B���/  �$�h��Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�2!  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �"  =�����.  �8A��`�E�;���  }�ع�B�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��K
3��E��EԉE؉E܋E΋��  3�#�#ʁ� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uB�E����u9u�u9u�u3�f�E���  f;�u!B�C���u9su93u�ủuȉu���  �u��}��E�   �E��M���M���~R�DĉE��C�E��E��M��	� �e� ���O��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?�����  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋M��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9M�w�Mԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�B�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�U�f�EċE؉EƋE܉E�f�U��3�f�����e� H%   � ���e� �Ẽ}� �<����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[�[���Ð:������\��������m�b����U���t�13ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�f��t�C-��C �u�}�f��u/��u+��u'3�f;�����$ f��C�C�C0�S3�@�  ��  f;���   3�@f��   �;�u��t��   @uhd�Qf��t��   �u��u;h\�;�u0��u,hT�CjP�Y�����3���tVVVVV�.������C�*hL�CjP�-�����3���tVVVVV�������C3��q  �ʋ�i�M  �������Ck�M��������3���f�M�8A�ۃ�`�E�f�U�u�}�M�����  }��B�ۃ�`�E�����  �E�T�˃������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE��P
3ɉM��M��M�M��M��3�� �  �u���  #�#֍4
����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��{����M�����?  ��  f;���  �E�3҉U��U��U�U��U��ɋ�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��V���3�3�f9u���H%   � ���E��\���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �^�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[��Q���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95�_��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��S  Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[�����U��SVWUj j h��u�  ]_^[��]ËL$�A   �   t2�D$�H�3��6M��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�d�5    �13�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�u�Q�R9Qu�   �SQ�`?�SQ�`?�L$�K�C�kUQPXY]Y[� ���������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ��U��j
j �u������]�������Q�L$+ȃ����Y��  Q�L$+ȃ����Y��  ��U��MS3�;�VW|[;�_sS������<� `�������@t5�8�t0�= Eu+�tItIuSj��Sj��Sj��� ���3���V���� 	   �^�������_^[]Ë�U��E���u�B����  �'���� 	   ���]�V3�;�|";�_s�ȃ����� `����@u$�����0����VVVVV� 	   �o���������� ^]�jh�$��v���}����������4� `�E�   3�9^u6j
�W���Y�]�9^uh�  �FP�����YY��u�]��F�E������0   9]�t���������� `�D8P�� �E��v���3ۋ}j
����YË�U��E�ȃ����� `���DP�� ]Ë�U����13ŉE�V3�95p?tO�=�C�u�"  ��C���u���  �pV�M�Qj�MQP���ug�=p?u�� ��xuω5p?VVj�E�Pj�EPV�P�� ��C���t�V�U�RP�E�PQ� ��t�f�E�M�3�^�;I�����p?   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��|T���E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�R���YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�� ���E�u�M;��   r 8^t���   8]��e����M��ap��Y����h���� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�� ���:���뺋�U��j �u�u�u�������]�����������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��jh�$��s��3ۉ]�j腍��Y�]�j_�}�;=�_}W������O�9tD� �@�tP�  Y���t�E��|(��O��� P�l ��O�4�*P��Y��O�G��E������	   �E��s���j�&���YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV����YP�p�����;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�L���P�  Y��Y��3�^]�jh�$�r��3��}�}�j�3���Y�}�3��u�;5�_��   ��O��98t^� �@�tVPV�Q���YY3�B�U���O���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��uࡠO�4�V�Z���YY��E������   �}�E�t�E��r���j蜊��Y�j����YË�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�.  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�  �EPSj �u��M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�5  Y����  �t�Etj�  Y����v  ����   �E��   j��  �EY�   #�tT=   t7=   t;�ub��M����D��{L�H��M�����{,�D�2��M�����z�D���M�����z� D�� D��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�  �M��]�� �����������}�E�����S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj�   Y�e���u��Et�E tj �   Y���3���^��[�Ë�U��}t~�}譄��� "   ]�蠄��� !   ]�3�Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-l@�]���t����-l@�]�������t
�-x@�]����t	�������؛�� t���]����jh%��k��3�9�_tV�E@tH9�@t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�@ �e��U�E�������e��U��k��Ë�U����13ŉE�j�E�Ph  �u�E� �� ��u����
�E�P�6���Y�M�3��)?���Ë�U���4�13ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5� �M�QP�֋� ��t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u�讥����YF;�~[�����wS�D6=   w/������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P��E��Y;�t	� ��  ���E���}�9}�t؍6PW�u��F����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�� ��t`�]��[�� 9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�\��YY�E�;�t+WWVPV�u�W�u��;�u�u��zF��Y�}���}��t�MЉ�u�����Y�E��e�_^[�M�3��u=���Ë�U����13ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[�;����3�PPjPjh   @ht���Cá�CV�5���t���tP�֡�C���t���tP��^Ë�U��SV�uW3����;�u�Q��WWWWW�    ��~������B�F�t7V�����V���M  V�о��P�t  ����}�����F;�t
P��C��Y�~�~��_^[]�jh(%��f���M��3��u3�;���;�u��~���    WWWWW�V~���������F@t�~�E���f���V�p���Y�}�V�*���Y�E��E������   �ՋuV辽��Y�jhH%�xf���E���u�^~��� 	   ����   3�;�|;�_r�=~��� 	   SSSSS��}�����Ћ����<� `��������L��t�P�8���Y�]���Dt1�u����YP���u� �E���]�9]�t��}���M��}��� 	   �M���E������	   �E���e����u�n���YË�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$�I������"Q���EQQ�$�4��������  �����  �E�]���������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U��V�uWV�����Y���tP� `��u	���   u��u�@Dtj�����j������YY;�tV����YP���u
� ���3�V���������� `����Y�D0 ��tW��{��Y����3�_^]�jhh%�c���E���u�{���  �{��� 	   ����   3�;�|;�_r!�w{���8�]{��� 	   WWWWW��z�����ɋ����� `��������L1��t�P�X���Y�}���D0t�u�����Y�E���{��� 	   �M���E������	   �E��6c����u����YË�U��V�u�F��t�t�v�?���f����3�Y��F�F^]�����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%� ������������h���^@��Y����̃=�D uK��D��t��D�Q<P�B�Ѓ���D    ��D��tV��萞��V躝������D    ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �& �&  ' ' ' .' :' L' `' t' �' �' �' �' �' �' ( ( ( 4( D( \( d( r( �( �( �( �( �( �( �( ) .) D) ^) l) z) �) �) �) �) �) �) * * .* <* H* T* ^* j* |* �* �* �* �* �* �* + + ,+ <+ N+ `+ p+ �+ �+ �+ �+ �+ �+         ��        �;.b����        ��5�                    �0N       p   � � bad allocation  USERNAME      zD         @�@ikto    ikfrom  texturesearchpath   dst src 
�#<fbx c4d EXPORT_ERROR: An unknown error has occured  EXPORT_ERROR: An error occured while saving the document    EXPORT_ERROR: Destination bad format    EXPORT_ERROR: Source bad format EXPORT_ERROR: Source either does not exist or cannot be located EXPORT_ERROR: An error occured while loading the document   EXPORT_ERROR: FBX exporter not found    SUCCESS framerate=  version=    -UnityC4DFBXtmp -UnityC4DFBXout 0   Filtered:       Name: ' '   Plugin:     Processing  Scanning    -UnityC4DFBXcmd * (c) 2006-2011 Unity Technologies ApS - http://unity3d.com * Unity-C4DToFBXConverter for Cinema 4D R11. Version: 3.09  ����MbP?l p� �f � P� %s      !@�  B   KB  MB       P? GB #   M_EDITOR    �������^          �?        O1\\    H!�7e+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    E`EEncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:    ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx                            �?5�h!���>@�������             ��      �@      �            	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        ������tl`T��|hH,LD(@<840,  ��������������������������x`T@  ���|`<��������tdH( ���hD ����GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                                                                                                                                                                                                                                                                                             ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun 1#QNAN  1#INF   1#IND   1#SNAN  _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   modf    fabs    floor   ceil    tan cos sin sqrt    atan2   atan    acos    asin    tanh    cosh    sinh    log10   log pow exp SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$     H                                                           1�!   RSDS��S�Y�E��	I�-   C:\BuildAgent\work\b2b44f52c74c2f2a\src\obj\Unity-C4DToFBXConverter11_Win32_Release.pdb            H P     l0        ����    @   8             �0�            � �     �0        ����    @   �             �0�            � � P     �0       ����    @   �             �0!           $!,!    �0        ����    @   !            41\!           l!t!    41        ����    @   \!�] d� �                     ����    ����    �����3�3    ����    ����    ����    �8    ����    ����    ����    �:    ����    ����    ����    "<    ����    ����    ����    KL����    ZL����    ����    ����    N����    N����    ����    ����    �S    ����    ����    ����OVSV    ����    ����    �����a�a    ����    ����    ����    �b    ����    ����    ����    ?w    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    y�    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    X�    ����    ����    ����[�o�    ����    ����    ��������    ����    ����    ����    ��    ����    ����    ����(�?�    ����    ����    ����    ��    ����    ����    ����    ǲ    ����    ����    ����    K�    ����    ����    ����    A�    ����    ����    ����    ��        ������    ����    ��������    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ���%         �&                        �& �&  ' ' ' .' :' L' `' t' �' �' �' �' �' �' ( ( ( 4( D( \( d( r( �( �( �( �( �( �( �( ) .) D) ^) l) z) �) �) �) �) �) �) * * .* <* H* T* ^* j* |* �* �* �* �* �* �* + + ,+ <+ N+ `+ p+ �+ �+ �+ �+ �+ �+     ZGetTempPathA  KERNEL32.dll  �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �GetLastError  �HeapFree   GetProcAddress  �GetModuleHandleA  -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent �GetModuleHandleW  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �InterlockedIncrement  �SetLastError  �InterlockedDecrement  !Sleep ExitProcess �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA � DeleteCriticalSection �GetModuleFileNameA  JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW zWideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy WVirtualFree TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �WriteFile �LeaveCriticalSection  � EnterCriticalSection  TVirtualAlloc  �HeapReAlloc �HeapSize  [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �LoadLibraryA  �InitializeCriticalSectionAndSpinCount �RtlUnwind �GetLocaleInfoA  �SetFilePointer  �GetConsoleCP  �GetConsoleMode  �LCMapStringA  MultiByteToWideChar �LCMapStringW  =GetStringTypeA  @GetStringTypeW  �SetStdHandle  �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW ZRaiseException  x CreateFileA C CloseHandle AFlushFileBuffers              �0N    ",          , ,  , �. @,   Unity-C4DToFBXConverter11.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                        |    |    B�     b�     a�     `�     ��    ��    qr            |||||||�    .?AVGeSortAndSearch@@   �    .?AVNeighbor@@  �    .?AVDisjointNgonMesh@@  |||||�    .?AVBaseData@@  |||||||||u�  s�  N�@���D            |�    .?AVtype_info@@     sqrt    �������������������S    �����
                                                                   x   
   |                  H   	   �

   X
   ,
   �	   �	   �	   t	   L	   	   �   �   �   0    �!    "   `x   Ly   <z   ,�   (�   ��                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                                  ���5�h!����?      �?                                                                                                                                                                                                                                                                                                                                          abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     �5�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����C                                                                                              �:            �:            �:            �:            �:                              �>        � (>�:   �:�5        �O    �O                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HD@<840(  ����������������������tl`TPL@, 	         (>.   �>�N�N�N�N�N�N�N�N�N�>   .                 ���5      @   �  �   ����              �                              0   ,   (          !          �   �   �   �   �   �    �   �   �   �   �   �   �   �   �   �"   �#   �$   �%   x&   l�&         �D        � 0     �p     ����    PST                                                             PDT                                                             �@�@����        ����                 �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
��������          �      ���������              �����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                                                                                                                                                                                                                                                                                                                                                                                     �   0"000A0N0d0�0�0�0�01191I1t1�1�1�1S2s2�2313G3�3�3�3�3�34%4F4S4b4j4�4�4�4�4�4r5�5�5�56/6�6�6�6�6�67*7N7�7�78)8W8�8�8949P9k9|9�9�9�9�9::1:C:m::�:�:�:�:�:�:;;.;N;\;t;�;�;�;�;�;<<.<N<h<�<�<�<�<�<�<==`=g=�=�=�=�=�=>->?>W>�>�>3?L?�?    (  0@0�0�0�0\12=2W2�2�2�2353G3Y3�3�3�3�3�3*4<4M4_4q4�4�4�4�45�5�5�56616E6Z6o6�6�6�6�6�6�6�67)7>7g7n7�7�7�7�7	8'8G8e88�8�8�8�8�8�8�899.9?9`9�9�9+:E:d:h:l:p:t:�:�:�:�:�: ;;;2;;;L;a;j;|;�;�;�;�;�;�;�;:<X<p<�<�<�<�<�<�<=^=s=�=�=�=�=�=�=>.>F>n>t>�>�>�>�>�>�>?*?@?Q?c?l?�?�?�?�?�?   0     00(010F0[0t0�0�0�0�0�0�0�01L1_1~1�1�1�1�1�1�1 24282<2@2D2H2L2P2T2X2\2`2�2�2�2�2�2�2�233(3r3�3�3�3�3�34#454G4Y4k4|4�4�4�4�455-5?5Q5c5t5�5�5�5�5�56 616Q6|6�6�6�67*7<7�7�7�7�7�7�788;8L8^8p8�8�8�8
9919H9Z9l9�9�9�9�9::%:7:H:�:�:�:�:;�;<2<e<�<�<=e=�=�=�=5>u>�>?O?�?�? @  �   0B0u0�01R1�1�12E2u2�2�2%3U3�3�354u4�4�45@5T5d5�5�56U6�6�6%7e7�7�7898C8m8r8�8�8�89)9e9�9�9�9E:i:�:�:�:&;O;�;�;�;<V<�<='=D=d=�=�=�=�=>>$>A>Q>d>�>�>�>�>�>?1?Q?t?�?�?�? P  �   0$0D0d0�0�0�011$1D1d1�1�1�1�122D2o2�2�2�23 3A3T3t3�3�3�3�3!4A4a4�4�4�45D5�5�56$6D6d6�6�6�6�6747T7�7�7�7�7'8D8q8�8�8�89A9d9�9�9�9!:t:�:�:�:4;T;t;�;�;�;<4<Q<t<�<�<�<=1=T=�=�=>!>D>d>�>�>�>?!?A?a?�?�?�? `  �   0$0T0q0�0�0�0D1�1�1�1242d2�2�2�2313Q3q3�3�3�3444d4�4�4�4$5[5�5�5�5�56D6t6�6�6�6�6
7$7t7�7�7�748T8�829�9�9�9
:-:a:�:�:�:;/;t;�;�;=$=Q=t=�=�=>>7>T>�>�>�>�>?4?d?�?�?�?�? p  �   10T0�0�0�0�0141q1�1�1�1D2�2�23!3D3d3�3�34a4~4�4�4�4525[5l5�5�5�5�5626Z6n6�6�6�67%7Z7m7�7�7�7�7�7�8�859V9�9�;�=�=�=B>�>�>�> �  �   <0@0D0H0{0�0�0�0�01D1d1�1�1�1�1242T2t2�2�2�2�2�2�2343T3t3�3�3�3444T4t4�4�4�4�4�45$5D5d5�5�5�5�5646Q6d6�6�6�6�67$7d7�7�7�7�7848T8t8�8�8�8�8949T9t9�9�94:c:�:�:4;a;�;�;�;<<D<d<�<�<�<�<�<=$=D=y=�=�=>%>H>t>�>�>�>?2?F?V?�?�?�?�?�?   �     040T0t0�0�0�0�0141i1}1�1�1�12222B2d2~2�2�2�23D3\3�3�3�3�34c4u4�4�4545T5t5�5�5�56$6D6d6�6�6�6�6�6$7D7d7�7�7�7	848T8t8�8�8�8�8	9959F9X9t9�9�9�9�9:%:D:U:t:�:�:�:�:�:$;Q;t;�;�;�;�;�;<<4<T<t<�<�<�<�<=D=d=�=�=�=>>4>a>t>�>�>�>?D?d?�?�?�?�? �  �   040T0t0�0�0�0�0141W1�1�1�1�1�12t2�2�2�2�243Q3�3�3�3�34+4$5D5d5�5�5�5�56$6Q6a6t6�6�6�6�6�6737A7P7q7�7�7�78!8A8Q8a8t8�8�8�8�8	9 9/9T9t9�9�9�9�9:4:T:t:�:�:�:�:�:;4;G;`;o;�;�;�;�;�;A<T<�<�<�<�<=4=T=t=�=�=�=�=>4>T>t>�>�>�>�>?4?d?�?�?�?   �  �   040T0t0�0�0�0�0$1D1t1�1�1�1�1242T2t2�2�2�23$3D3d3�3�3�34!4A4d4�4�4�4�4�4545I5`5o5�5�5�5�5646d6�6�6�67T7x7�7�8�8�8�8�89o9�9�9�9::1:M:x:�:�:�:�:;!;D;d;�;�;�;�;<$<T<�<�<�<=$=Q=a=�=�=�=�=>$>I>d>�>�>�>�>$?N?t?�?�?�?�?   �  �   0D0�0�0�041U1f1�1�1�1�1�1�1�1$2^2�2�2�243T3�3�3�3444k4�4�4�4�4545T5t5�5�5�5$6D6Z6�6�6�67D7t7�7�7�7818Q8d8�8�8�8�8$9?9_9r9�9�9�9�92:T:t:�:�:�:�:;4;d;�;�;�;<$<d<�<�<�<=$=D=d=�=�=�=�=>!>4>T>t>�>�>?>?S?�?�? �  �   Q0w0�0H1j1�12*2M2�2�2�2n3�3�3#4L4i4�4�4�4�5�5�5C6l6�67,7I7�7�7�7k8�89a9�9�9:a:�:�:L;�;�;	<~<�<�<.=N=c=�=>|>�>?4?Q?a?t?�?�?�?   �  �    0$0T0t0�0�01$1D1a1�1�1�1C2`2�2�2�2�2	3F3U3�3�3�3�3444�4�4�4�4�4!5D5d5�5�5�5�5646d6�6�6�67!777|7�7�78\8�8�8�89!919D9�9�9�9�9�9:$:L::�:&;E;�;�;)<E<�<�<-=E=�=>5>�>�>,?H?l?�?�?�?�?   �  D  0,0H0l0�0�0�0�01$111_1�1�1�1�12,2\2�2�2�2�2�2343J3x3�3�3�3 4Q4c4u4�4�4�4�4#5C5W5o5�5�5�5%6d6�6�67)7T7]7j7�7�7�7�7�7�7�7�78%8B8T8p8�8�8�8�8�8�8�89)9;9M9_9h9�9�9�9�9�9::%:.:J:g:x:�:�:�:�:�:;";/;G;Y;k;};�;�;�;�;�; <<2<C<U<^<z<�<�<�<�<�<=="=>=\=n=�=�=�=�=>>'>9>K>]>o>x>�>�>�>�>�>?#?5?>?Z?w?�?�?�?�?�?�?     |   00<0N0j0�0�0�0�0�01-1T1q1�12
22&202K2g2�2�2�2�2�23F3l3�384M4p4�4�5�5�5�56$6D6d6�6�6�6�6747T7q7�7�7�78�8�8    $   �1�1�214f495o5�5�>�>?E?�?�?   t   0U0�0�0151u1�1�1%2e2�2�23B3r3�3�3%4u4�45E5�5�56e6;x;|;�;�;�;�<-=�>�>�>�>�>?!?;?o?�?�?�?�?�?�?�?�?�?�? 0 �   010_0�0�0�0�0�0�01	11111"1(1,12161<1@1F1J1c1t1�1�1�1�122"2h2n2�2�2�2�2@3m3�3/4H4O4W4\4`4d4�4�4�4�4�4�4�4�4�4�4�4>5D5H5L5P5�5�5�5�5�5�5�56;6m6t6x6|6�6�6�6�6�6�6�6�6�6�6B7^7�7�8�899?9v9�9�9M:_:�:�:�:;;�;�;�;�;�;�<�<�<�<�<$=,=A=L= @    0s0�06�6d8�8�8�8�8�8�89!9'9-93999@9G9N9U9\9c9j9r9z9�9�9�9�9�9�9�9�9�9�9�9�9�9�9:::#:.:::O:V:j:q:�:�:�:�:�:�:�:�:;;;";1;7;@;L;Z;`;l;r;;�;�;�;�;�;�;�;<)<i<o<�<�<�<�<�<s=�=�=�=�=,><>B>N>T>d>j>>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????"?(?,?2?7?=?B?Q?g?r?w?�?�?�?�?�?�?�?�?�?�? P   0:0C0O0�0�0�0�0�0�011C1^1d1m1t1�1�1�122 202:2A2L2U2k2v2�2�2�2�2�2	33@3E3P3U3s3�344)4J4P4�4�4�4!5+5S5l5�5�5�5A6G6k6�6�6�6�6�67W7b7l7}7�7;9L9T9Z9_9e9�9�9�9�9::(:/:f:�:�:�:;";';H;M;�;�;�;�;�;�;�;�;�;�;�;�;�;<<*<�<�<�<�<�=�=>�>�>�>?k?�?�?�?�?�?�?�? ` `   0	0142>2^2c2D3O3r364C4f4�4�4�4�4�4�4�4=5B5j5�5�5�5�5�56<6F7M7X8�89>9�9�9�9=>�?�?�? p �   �1�3�3�3�3�3�3�3�3�3�3�4�4�45
5"5N5j5�5�5�5�5�566"6E6L6e6y66�6�6�6T7t7�7�7�9�9�9�9�9::":-:?:R:]:c:i:n:w:�:�:�:�:�:�:�:�:�:�:�:�:�:;;; ;:;K;Q;b;�;c?o?�?�?   � �   0G02%2-2H2U2_3�3�3�3)4�485�5k6l7|7�7�7�7�7O8�8�8:':a:n:x:�:�:�:�:�:�:�:;;<;s;�;�;+<H<�<�<=�=�=�=�=�=�=�=>>8>A>G>P>U>d>�>�>�>�>�?�?   � �   "0n0�01k1�1�1�1M2Y2�3�3f4:5o5�5�5�5�5�5�5�5�5666 6$6(6,60646~6�6�6�6�6�677#7(7,707Q7{7�7�7�7�7�7�7�7�7�78 8$8(8,8�:�<�<[=p=�=�=�=>P>�>�>�>J?P?t?�?�?�?�? � �   $0�0�0�01!1'1�1�1�1�1�1�1�1�1.2<2�2�2�2�2�2�2�2�2Y3b3h3�34
44O4�4�46=6K6Q6a6f6~6�6�6�6�6�6�6�6�6�6�6�617N7k7�8�8�8h9u9�9�9�9:�:7;�;<�<$=}=?�? � �   �0�0�0<1[1�1,2[2�2?3l33�3�3�3�3�3�3�3�3�34*4<4J4_4i4�4�4�4�4�4-5f5q5�6�6':.:]:Q;�;�;�;�;�;�;�;�;/<�<v=�=>�>p?z?�?�?�?�?�?�?�? � T   �0�0
33.3P3b3t3�3�3�3�3�5�6�6E7'8�8�8h9n9~9:5:�:�;�;�<k=>
>�>�>�>b?y?�?   � 4   6033h6l6p6t6x6|6�6�6�6�6�6�6�6|7�7�7�7/8S8 � p   ]24m4y4�455�5�5�56p6�6�6�637>7l7z7�7�7�7�7�7�7�7�7�78
8 8;8�8N9�9�9�9:::":�: ;+;N;�;>i?�?�?�?�? � `   #0I1[1m1�1�1�1�12(2T2�2�2y3�34�5�5�5�5�56�67;7c7�7�7X9�9�9�9�9:C:�;�;�;�;�;�; <<     4   $1014181<1H1L1H4L4P4T4X4d4h4�4�4�4�4�455    �   �2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4�?�?   �   D0H0P0h0x0|0�0�0�0�0�0�0�0�0�0�0�011 1$1,1D1T1X1h1l1t1�1�1�1�12(2H2T2p2|2�2�2�2�2�2�2383X3x3�3�3�3�3�34484T4X4x4�4�4�4�455 5@5`5�5   0 @   00P0T0X0\0`0d0h0l0�0�0�0�0�0�0�0�0�0�0�0�0 111110141X1\1`1d1h1l1p1t1x1|1�1�1�12222$2,242<2D2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�9�:;;(;8;H;l;x;|;�;�;�;�;�;�;�; >$>(>,>0>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ?????�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? @ (   0000$0,040<0D0L0T0\0d011                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  