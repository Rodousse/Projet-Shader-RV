MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �	Q��h?�h?�h?�'��h?���h?����h?艮D�h?�h>��h?���h?���h?���h?�Rich�h?�                        PE  L 9	0N        � !	  
  �      �8                               �                               O Y   �H (                            � �  `!                            �B @                                         .text   	     
                   `.rdata  y/      0                @  @.data   �2   P     >             @  �.reloc  �&   �  (   V             @  B                                                                                                                                                                                                                                                                                                                                                                                        U��E��dt���   uB�`f    ]áhf�H�Q4��+`f=�  |�0(  �hf�H�Q4�ң`f�   ]��������U��hf�UV��H�AVR�Ѓ���^]� ��������������U��hfV��H�QV�ҡhf�H�U�AVR�Ѓ���^]� U��hfV��H�QV�ҡhf�U�H�E�IRj�PV�у���^]� ����������U��hf�P�E�RP��VWP�EP�E�P�ҋu���hf�H�QV�ҡhf�H�QVW�ҡhf�H�A�U�R�Ѓ�_��^��]� ���������������U��hf�P�R`��VW�E�P�ҋu���hf�H�QV�ҡhf�H�QVW�ҡhf�H�A�U�R�Ѓ�_��^��]� �������U��hf�H�U�I(��VWR�E�P�ыhf�u���B�HV�ыhf�B�HVW�ыhf�B�P�M�Q�҃�_��^��]���U���8�EV�]�W�E3��]�3��E �]��3��U���  �E�E�M�E�P�M�Q�M��E�   �U��E�   �9  �U�R��� >  ����u�E�PS�D  ��������   V���;>  �hf���   ���   jj���Ћ���tX�hf���   �E�Rlj P���҅�t;�hf�D�ȋ��   ���$�ȋB0V�ЍM��X*  G���.���_�   ^��]ÍM��;*  _3�^��]����U��QV�u���QO  �E���t}���$    ��hf���   �ȋB��=/  t)-�  t"���=��t�hf���   �M��B(���'�hf���   �M��BL�ЍM�Q�F  ������N  �E���u�^��]���������U��V�u��tB��I V�J����hf���   �B4������P������hf���   �B(�����Ћ���u�^]�U��hf�H�A�� S�U�VR�Ћhf�Q�J�E�P�ыhf�B�Pj j��M�h�!Q�ҍE�P�M�Q�݌  �hf���B�P�M�Q���ҋu��$V��t@�hf�H�Q�ҡhf�H�Qj j�h�!V�ҡhf�H�A�U�R�Ѓ���^[��]Ëhf�Q�B�Ћhf�Q�J�E�VP�ыhf�B�P�M�Q�҃���^[��]��������������U���0  � Q3ŉE�V�u��袏  ������Ph  �  ��t������Q������誏  �������jR誤  ��P����  �������D�  �M���3�^��  ��]����U��Q����L  �E�����   ���$    ��hf���   �ȋB�Ћhf=L  uN�Q@�E��J,P�у�h�  ���E�  ��u)�hf���   �M��PL�ҍE�P�4D  �����jL  ��hf���   �M��B(�ЉE����y�����]������U��V�u��t>��I �;����hf���   �B4����P������hf���   �B(�����Ћ���u�3�^]�����  P����Y����U���`SV�uW����  �}�]��    ����  �hf���   �Bx���Ћhf���   �E�Bx���Ћhf�Q�M�RxQ���҅��w  �hf���   �B����=  ��   �hf���   �B����=  ��   �hf�QH�R`�E�P����� �]���@�]��@�hf�PH�]��Rp�E�P��� �]Ћ��@�]��@�hf�PH�]��Rh�E�P��� �]����@�]��@���]�h�  �E�W��E��X�E��X�;����EЃ����h�  �E�W�X�E��X�����E������h�  �E�W�X�E��X������� �hf���   �B4���ЋM�UWQRP�hf���   �B4����P�R����hf���   �B(�����Ћhf���   ���B(���Ћ؅��=���_^[��]�������U����hf���   �SVW�}j j �������]������]���  P������]��;]�]�E���]��K�  �E�E���M��}���!�����]��$�w�  �M�Q���,�  �U�R���!�  j jjjj ����  �E�PVW���s�  P���k�  P�U���C��;]�]~�����]�M���!�$��  �M�Q�����  _��^[��]�������������U��hf�P�B<��D�M�Ѕ�u�hf�Q�J�EP�у�3���]Ëhf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q���   ��j �E�Pj=�M�҅�u>�hf�H�A�U�R�Ћhf�Q�J�E�P�ыhf�B�P�MQ�҃�3���]ËM�V�E�PQj �U�R�M������������hf�Q�R�M�QP�ҡhf�H�A�U�R�Ћhf�Q�J�E�P�ыhf�B�P<���M�ҋM�+�HPAQ�E�P�M�����hf�Q�R�M�QP�ҡhf�H�A�U�R�Ћhf�Q�E�RP�M�Q�ҡhf�H�A�U�R�Ћhf�Qj j�h�!�E�P�J�ыhf�B�Px��(�M�Q�M��ҋ�hf�H�A�ލU��RF�Ѓ���tB�hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�A�UR�Ѓ��   ^��]�j h�!�M�������hf�Q�Rx�E�P�M��ҋ�hf�H�A�ލU��RF�Ѓ���tB�hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�A�UR�Ѓ��   ^��]�j h�!�M��g����hf�Q�Rx�E�P�M��ҋ�hf�H�A�ލU��RF�Ѓ���tB�hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�A�UR�Ѓ��   ^��]�j h�!�M�������M�Q�M��  �hf���B�P�M�Q�҃���tB�hf�H�A�U�R�Ћhf�Q�J�E�P�ыhf�B�P�MQ�҃��   ^��]�j h�!�M��j����E�P�M��  �hf�Q�J���E�P�ыhf�B�P�M܃�Q�ҡhf�H�A�U�R�Ћhf�Q�J�EP�у���t
�   ^��]�3�^��]�����������U���tSV3�W95Pt)�P�jS�~�  ������uBF9<�P��Pu܍M�̇  �M$�ć  �hf�Q�J�E@P�у�_^�'  [��]Å�tˍEj P��  ����u1�M腇  �M$�}�  �hf�Q�J�E@P�у�_^�'  [��]Ëhf�B�P�M�Q�ҡhf�H�A3�Vj��U�h�!R�Ѓ��M�Q�M���  �hf���B�P�M�Q�E��҃��}� �Mt-���  �M$��  �hf�H�A�U@R�Ѓ�_^�'  [��]�VjQ�u��S�  ���E��M;�u.豆  �M$詆  �hf�B�P�M@Q�҃�_^�'  [��]ÍE�P过  �M�P�6�  �M��n�  �M$��  ���  �M$Q�M肆  �M$�ڈ  Vh�!�M������U�R�M$���  �hf�H�A�U�R�Ѓ��M$VQ蒕  ����t�U$VR���  ���M���  P�p����M����U�  �Mģdf�X�  �hf�E�    ���   �R�E�Pj���ҋE���>  �hf�Q@P�B,�Ћ������"  �hf�Q���   j j �E�P���ҡhf�P�B0jh�  ���Ћhf�Q�B0jh�  ���Ћhf�Q�B0j h�  ���Ћhf�Q�B0jh�  ���Ћhf�Q�B0j h�  ���Ћhf�Q�MP�R03�;MT����Ph�  ���   Vh�!�M������M�Q�M$蕇  �hf���B�P�M�Q�E��҃��}� ������M蘄  �M$萄  �hf�H�A�U@R�Ѓ�_^�'  [��]ËEP�MT;�}QP�E�P�+������E��M�j	Q�
n  �U�jR��m  ���E�P�M�p�  Pj	�n  ���M���  �hf�Q�B<�M@�Ѕ�t"�M@Q�M��|�  �U�Rj��m  ���M���  �M�Sj �E$PQ���  ������t�hf�B���   j j V�M��ҍE�Pj	�m  �M�Qj�m  �U�R�վ  ���M�芃  �M�肃  �M��Z�  �M�r�  �M$�j�  �hf�H�A�U@R�Ѓ������_%����^'  [��]����������������U����  ��  �E��E�P�f����� ���Q�Z����hf�B�P<���M��҅���  �hf�H�A�U�R�Ћhf�Q�Jj j��E�h�#P�эU�R�E�P�M�Q�a  �� P�M��%�  P�� ���R�����P��  ���M�膂  �hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h�#P�эU�R�E�P�M�Q��  ��(P�M�虁  P�� ���R������P�e�  ���M����  �hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h�!P�ыE��='  ��  ��  ����  WPh�#��,����Y���j h�#������G���j h|#��<����5����hf�:�EP�M�Q�g  ��P������WR������P��,���P������Q�hg  �df��PR������P�������P�����Q��D���R�:g  P��<���P������Q�  ��P��$���R�v  ��P������P�f  ��P��d���Q�V  ��P��4���R�F  ��P��T���P�6  ��P��t���Q�&  ��P������R�  ��P�M�������hf�H�A������R�Ћhf�Q�J��t���P�ыhf�B�P��T���Q�ҡhf�H�A��4���R�Ћhf�Q�J��d���P�ыhf�B�P������Q�ҡhf�H�A��$���R�Ћhf�Q�J������P�ыhf�B�P��D���Q�ҡhf�H�A������R�Ћhf�Q�J������P�ыhf�B������Q�P�ҡhf�H�A�U�R�Ћhf�Q�J��<���P�ыhf�B�P�����Q�ҡhf�H�A��,���R�Ѓ�@_��  j hT#�M�������hf�Q�R�E�P�M�Q�ҡhf�H�A�U�R�Ѓ��  �������0  �$�$* j h#��\���������\���Q�M������hf�B�P��\���Q�҃��A  j h�"��L����G�����L���P�M�������hf�Q�J��L���P�у��  j h�"��l����	�����l���R�M������hf�H�A��l���R�Ѓ���   j h�"��|����������|���Q�M��]����hf�B�P��|���Q�҃��   j hT"�M������E�P�M��%����hf�Q�J�E�P�у��V�hf�B�P�M�Q�ҡhf�H�Aj j��U�h("R�Ћhf�Q�R�E�P�M�Q�ҡhf�H�A�U�R�Ѓ� �hf�Q�J�E�P�ыhf�B�Pj j��M�h�!Q�ҡhf�H�I�UR�E�P�ыhf�B�P�M�Q�ҡhf�E�    �H���   h�!h�   h   �ҋhf��,j �E��Qh   P�Bh�M���h1D4ChCD4Cjj j������Q�M�萁  �hf�B�Pdj �M��ҋM�P�E�P���  �M�舁  j�����Q������R�#�  ������j P���  �M�Q���  �hf�B�P�M�Q�҃��������|  ������|  �� �����{  �hf�H�A�U�R�ЍM�Q輀  �hf�E�    �B�P�MQ�҃���]�)' g' �' �'  ( ��������U����   SVW�_�  h1D4ChCD4Cjj j�MQ�ȉE�聀  �hf�B�P�M�Q�ҡhf�H�Aj j��U�h�!R�Ћhf�Q�J�E�P�ыhf�B�Pj j��M�h�!Q�ҡhf�H�A��x���R�Ћhf�Q�Jj j���x���h�!P�ыhf�B�P�M�Q�ҡhf�H�A��@j j��U�h�!R�Ћhf�Q�J�E�P�ыhf�B�Pj j��M�h�!Q�ҡhf�E� �H�A�U�R�Ћhf�Q�Jj j��E�h�!P�ыhf�B�P�M�Q�ҡhf�H�Aj j��U�h�!R�ЋM���L3���  ����  ����  3�3�j j�M�Q�M��[  �E�<
�4  <�,  �M���  ���� ;���  ;���  f�U��hf�H�A��8���R�Ћhf�Q�JV��8���jP�ыhf�B�P<���M��ҋhf�Q�RLj�j���8���QP�M��ҡhf�H�A��8���R�Ћhf�B���M�Q�H����V�ыhf�B�P�M�VQ�҃����������wq�$�42 j h�!���������������P�M��k����hf�Q�J�����P�у��/�U�R�M��!�M���M�Q��x�����U�R�M���M��E�P�"����hf�Q�J��X���P�ыhf�B�Pj j���X���h�!Q�ҡhf�H�I�U�R��X���P�ыhf�B�P��X���Q����  f�E��hf�Q�J����(���P�ыhf�B�PV��(���jQ�ҡhf�P�B<���M��Ћhf�Q�RLj�j���(���QP�M��ҡhf�H�A��(���R�Ѓ��j  �hf�B�M�Q�H����V�ыhf�B�P�M�VQ�҃��Y���������   �$�L2 �hf�H�A��H���R�Ћhf�Q�Jj j���H���h�!P�ыhf�B�@�M�Q��H���R�Ћhf�Q�J��H���P�у� �h�hf�B�@�M�Q�U�R���M�E��5�hf�H�I��x���R�E�P���.�hf�B�@�M�Q�U�R����E��hf�Q�RP�M�Q�҃��hf�H�A�U�R�Ћhf�Q�Jj j��E�h�!P�ыhf�B�@�M�Q�U�R�Ћhf�Q�J�E�P�у� �M�C�Ù�����2|  ;��/���;��%����M��X{  �Uj R�݅  �hf�H�A��h���R�Ћhf�Q�Jj j���h���h�!P�ыhf�B�P<���M��҅�uW�hf�H�A�U�R�Ћhf�Q�Jj j��E�h�#P�ыhf�B�@�M�Q�U�R�Ћhf�Q�J�E�P�у� �hf�B�P<�M��҅�uW�hf�H�A�U�R�Ћhf�Q�Jj j��E�h�#P�ыhf�B�@�M�Q�U�R�Ћhf�Q�J�E�P�у� �hf�B�PXj �M��ҋ�hf�P�BXj �M��Ћhf��h���QVP�B�H����V�ыhf�B�P��x���VQ�҃��E���P�(t  ���U���R�t  �������hf�H�Q��D��V�ҡhf�H�A��h���VR�Ѓ�W�2����hf�Q�J��h���P�ыhf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q�E��JP�ыhf�B�P�M�Q�ҡhf�H�A��x���R�Ћhf�Q�J�E�P�ыhf�B�P�M�Q�ҍE�P�x  ��8�M�E�    �s  _^[��]��, - - - )- 2- j. �. �. �. / / ������������U���   SVW�/�  �����p  ��I �hf�H�A�U�R�Ћhf�Q�Jj j��E�h�#P�эU�R�[  �hf�H�A�U�R�Ћhf�Q�J�E�P�ыhf�B�Pj j��M�h�#Q�ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h�#P�у�D�U�R��`���P���ܺ  ���Us  �hf�Q�J���E�P�ыhf�B�@�M�Q�U�R�Ћhf�Q���B<�M��Ћhf�Qj�j�WP�BL�M��Ћhf�Q�J�E�P�ыhf�B�@�M�Q�U�R�Ћhf�Q�B<���M��Ћhf�Q�RLj�j��M�QP�M��ҍE�P��Y  �hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q�J�E�P�у���`����q  �hf�B�P�M�Q�҃�����  �hf�Q�J(P��|���P�ыhf���B�P�M�Q�ҡhf�H�A�U�RW�Ћhf�Q�J��|���P�эU�R�Y  �hf�H�A�U�R�Ћhf���   �B(�� ���Ћ���������hf�Q�J�E�P�ыhf�B�Pj j��M�h�#Q�ҍE�P�X  �hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�Aj j��U�h�#R�ЍM�Q�XX  �hf�B�P�M�Q�ҡhf���   ���   ��j��jS��  ��D����  �hf���   ���   ��3��Ѕ���  �hf���   ���   V���Ћhf�Q�J���E�P�ыhf�B�Pj j��M�h�#Q�ҍE�P�W  �hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�Aj j��U�h�#R�Ћhf�Q�J�E�P�ыhf�B�Pj j��M�h�#Q�҃�D��|���P��`���Q���{�  ����o  �hf�E��B�P�M�Q�ҡhf�H�U�R�I�E�P�ыhf�B�P<���M��ҋhf�Q�M��RLj�j�QP�M��ҡhf�H�A�U�R�Ћhf�Q�R�E�P�M�Q�ҡhf�P�B<���M��Ћhf�Q�RLj�j��M�QP�M��ҍE�P�oV  �hf�Q�J�E�P�ыhf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q�J��|���P�у���`����'n  �hf�B�P�M�Q�҃���苶  �hf�Q�J(P�E�P�ыhf���B�P�M�Q�ҡhf�H�A�U�RW�Ћhf�Q�J�E�P�эU�R�U  �hf�H�A�U�R�Ћhf���   ���   �� ��F��;��w���_^[��]��������������U��E���   P�����M�Q�����hf�B�P<���M��҅�u"�M��5m  �hf�H�A�U�R�Ѓ�3���]Ëhf�Q�J�E�P�ыhf�B�Pj j��M�h $Q�ҍE�P�M�Q�U�R�  �� P��|����Nl  P�E�P�M�Q� p  ����|����l  �hf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q�J�E�P�ыhf�B�Pj j��M�h�#Q�҃��E�P�M��m  P�M�Q�U�R��   P�/T  �hf�H�A�U�R�Ћhf�Q�J�E�P�ыhf�B�P�M�Q�ҍE�j P�{  ��$��tZ�hf�B�P�M�Q�ҡhf�H�Aj j��U�h�#R�ЍM�Q�S  �hf�B�P�M�Q�ҍE���P�fk  �������M��k  �M��k  �hf�Q�J�E�P�у�3���]����U��hf�P�E�RxP�����@]� ���U��hf�H�QV�uV�ҡhf�H�U�AVR�Ћhf�Q�B<�����Ћhf�Q�M�RLj�j�QP���ҋ�^]��������̡hf� 8����W  ;��@����������U��hf���8�������W  v3���]Ë@�P�M�Q�ҡhf�H�Aj j��U�hL$R�ЍM�Q�pR  �hf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h$P�эU�R�)R  �hf�H�A�U�R�Ѓ�8�   ��]�����������������������������U��hf� 8���=W  v3�]ËE�� t��t-Vu�u��]����   ]ù�f���  �����]�����U��E�hf� ]��hlfPhD � �  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��hlfjhD �L�  ����t
�@��t]��3�]��������Vhlfj\hD ����  ����t�@\��tV�Ѓ���^�����Vhlfj`hD �����  ����t�@`��tV�Ѓ�^�������U��VhlfjdhD ����  ����t�@d��t
�MQV�Ѓ�^]� ������������U��VhlfjhhD ���y�  ����t�@h��t
�MQV�Ѓ�^]� ������������VhlfjlhD ���<�  ����t�@l��tV�Ѓ�^�������U��Vhlfh�   hD ����  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vhlfh�   hD ����  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��VhlfjphD ���i�  ����t�@p��t�MQV�Ѓ�^]� �pf^]� ��U��VhlfjxhD ���)�  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vhlfj|hD �����  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vhlfj|hD ����  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� �������������U���Vhlfh�   hD ���S�  ����t=���   ��t3�MQ�U�VR��hlfj`hD �&�  ����t�@`��t	�M�Q�Ѓ���^��]� �����̋���������������hlfjhD ���  ����t	�@��t��3��������������U��V�u�> t+hlfjhD ��  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0hlfjhD �a�  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��VhlfjhD ����  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��VhlfjhD �����  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vhlfj hD ����  ����t�@ ��tV�Ѓ�^�3�^���Vhlfj$hD ���l�  ����t�@$��tV�Ѓ�^�3�^���U��Vhlfj(hD ���9�  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vhlfj,hD �����  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vhlfj(hD ����  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vhlfj4hD ���\�  ����t�@4��tV�Ѓ�^�3�^���U��Vhlfj8hD ���)�  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vhlfj<hD �����  ����t�@<��t
�MQV�Ѓ�^]� ������������VhlfjDhD ����  ����t�@D��tV�Ѓ�^�3�^���U��VhlfjHhD ���i�  ����t�M�PHQV�҃�^]� U��VhlfjLhD ���9�  ����u^]� �M�PLQV�҃�^]� �����������U��VhlfjPhD �����  ����u^]� �M�U�@PQRV�Ѓ�^]� �������VhlfjThD ����  ����u^Ë@TV�Ѓ�^���������U��VhlfjXhD ����  ����t�M�PXQV�҃�^]� U��Vhlfh�   hD ���V�  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vhlfh�   hD ����  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vhlfh�   hD ����  ����u^]� �M���   QV�҃�^]� �����U��Vhlfh�   hD ���v�  ����u^]� �M���   QV�҃�^]� �����U��Vhlfh�   hD ���6�  ����u^]� �M���   QV�҃�^]� �����U��Vhlfh�   hD �����  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vhlfh�   hD ��  ����u�hf�H�u�QV�҃���^��]ËM���   WQ�U�R�Ћhf�Q�u���BV�Ћhf�Q�BVW�Ћhf�Q�J�E�P�у�_��^��]��U��Vhlfh�   hD ���&�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vhlfh�   hD ���ֿ  ����t���   ��t�MQ����^]� 3�^]� �U��Vhlfh�   hD ��薿  ����t���   ��t�MQ����^]� 3�^]� �U��Vhlfh�   hD ���V�  ����t���   ��t�MQ����^]� 3�^]� �Vhlfh�   hD ����  ����t���   ��t��^��3�^����������������U��Vhlfh�   hD ���־  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vhlfh�   hD ��膾  ����t���   ��t�MQ����^]� ��������U��Vhlfh�   hD ���F�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vhlfh�   hD �����  ����t���   ��t��^��3�^����������������VW��3����$    �hlfjphD 诽  ����t�@p��t	VW�Ѓ���pf�8 tF��_��^�������U��SW��3�V��    hlfjphD �_�  ����t�@p��t	WS�Ѓ���pf�8 tqhlfjphD �-�  ����t�@p��t�MWQ�Ѓ�����pfhlfjphD ���  ����t�@p��t	WS�Ѓ���pfV���������tG�]����E^��t�8��~=hlfjphD 讼  ����t�@p��t	WS�Ѓ���pf�8 u_�   []� _3�[]� ����������U��Vhlfj\hD ���Y�  ����t3�@\��t,V��hlfjxhD �7�  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vhlfj\hD �����  ����t3�@\��t,V��hlfjdhD �׻  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vhlfj\hD ��薻  ����tG�@\��t@V�ЋEhlfjdhD �E��E�    �E�    �`�  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vhlfj\hD ����  ����t\�@\��tUV��hlfjdhD ���  ����t�@d��t
�MQV�Ѓ�hlfjhhD �κ  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vhlfj\hD ��艺  ������   �@\��t~V��hlfjdhD �c�  ����t�@d��t
�MQV�Ѓ�hlfjhhD �:�  ����t�@h��t
�URV�Ѓ�hlfjhhD ��  ����t�@h��t
�MQV�Ѓ���^]� ��U���VhlfjthD ���ֹ  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���hlfj`hD 螹  ����t(�@`��t!�M�Q�Ѓ���^��]� �uhpf���_�����^��]� ������U���Vhlfh�   hD �E�  ����tU���   ��tK�M�UQR�M�Q�Ћu��P������hlfj`hD ��  ����t%�@`��t�U�R�Ѓ���^��]ËE�uP���k�����^��]�����U���Vhlfh�   hD ��賸  ����tR���   ��tH�MQ�U�R���ЋuP������hlfj`hD �z�  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    �'�����^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t�hf���   P�B@��]� �E��t�hf���   P�BD��]� �hf���   R�PD��]� �����U��hf�P@�Rd]�����������������U��hf�P@�Rh]�����������������U��hf�P@�Rl]�����������������U��hf�P@�Rp]�����������������U��hf���   ���   ]�����������U��hf���   ���   ]����������̡hf�P@�Bt����̡hf�P@�Bx�����U��hf�P@�R|]����������������̡hf�P@���   ��hf���   �Bt��U��hf�P@���   ]�������������̡hf�P@���   ��U��hf�P@���   ]��������������U��hf�P@���   ]��������������U��hf�P@���   ]��������������U��hf�P@���   ]��������������U��hf�P@���   ]��������������U��hf�P@���   ]��������������U��hfV��H@�QV�ҋM����t��#����hf�Q@P�BV�Ѓ�^]� �̡hf�PH���   Q�Ѓ�������������U��hf�P@�EPQ�JL�у�]� ���̡hf�P@�BHQ�Ѓ����������������U��hf�P@�EP�EP�EPQ�J�у�]� ������������U��hf�P@�EPQ�J�у�]� ����U��hf�P@�EP�EPQ�J�у�]� U��hf�P@�EPQ�J �у�]� ����U��hf���   �R]��������������U��hf���   �R]��������������U��hf���   �R ]��������������U��hf���   ���   ]�����������U��hf���   ��D  ]�����������U��hf�E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U��hf���   ���   ]����������̡hf���   �B$��hf�H@�Q0�����U��hf�H@�A4j�URj �Ѓ�]����U��hf�H@�A4j�URh   @�Ѓ�]�U��hf�H@�U�E�I4RPj �у�]�̡hf�H|�������U��V�u���t�hf�Q|P�B�Ѓ��    ^]��������̡hf�H|�Q �����U��V�u���t�hf�Q|P�B(�Ѓ��    ^]��������̡hf�H@�Q0�����U��V�u���t�hf�Q@P�B�Ѓ��    ^]���������U��hf�H@���   ]��������������U��V�u���t�hf�Q@P�B�Ѓ��    ^]��������̡hf�PH���   Q�Ѓ�������������U��hf�PH�EPQ��d  �у�]� �U��hf�H �IH]�����������������U��}qF uHV�u��t?�hf���   �BDW�}W���Ћhf�Q@�B,W�Ћhf�Q�M�Rp��VQ����_^]����������̡hf�P@�BT�����U��hf�P@�RX]�����������������U��hf�P@�R\]����������������̡hf�P@�B`�����U��hf�H��T  ]��������������U��hf�H@�U�A,SVWR�Ћhf�Q@�J,���EP�ыhf�Z��h��hE  �΋��q  Ph��hE  ���q  P��T  �Ѓ�_^[]����U��hf���   ���   ]�����������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�PL�E��  PQ�MQ�҃�]� ������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�BQ�Ѓ����������������U��hf�PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U��hf�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��hf�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��hf�PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U��hf�PX�EPQ�J�у�]� ����U��hf�PX�EPQ�J�у�]� ����U��hf�PX�EPQ�J�у�]� ����U��hf�PX�EPQ�J�у�]� ����U��hf�PX�EPQ�J$�у�]� ����U��hf�PX�EPQ�J �у�]� ����U��hf�PD�EP�EPQ�J�у�]� U��hf�HD�U�j R�Ѓ�]�������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�HD�	]��U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�HD�U�j R�Ѓ�]�������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�U�HD�Rh2  �Ѓ�]����U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�U�HD�RhO  �Ѓ�]����U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�U�HD�Rh'  �Ѓ�]����U��hf�H@�AV�u�R�Ѓ��    ^]�������������̡hf�HD�j h�  �҃�����������U��hf�H@�AV�u�R�Ѓ��    ^]�������������̡hf�HD�j h:  �҃�����������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E��hf���   �R�E�Pj�����#E���]�̡hf�HD�j h�F �҃�����������U��hf�H@�AV�u�R�Ѓ��    ^]�������������̡hf�HD�j h�_ �҃�����������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E��hf�E�    ���   �R�E�Pj������؋�]� ̡hf�PD�B$Q�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ���������������̡hf�PD�B(Q�Ѓ���������������̡hf�PD�BQ�Ѓ����������������U��hf�E�PH�B���$Q�Ѓ�]� ���������������U��hf�PH�EPQ���   �у�]� �U��hf�PH�EPQ���  �у�]� �U��hf�PH�EPQ���  �у�]� �U��hf�PH�EP�EPQ��  �у�]� �������������U��hf�PH�EP�EPQ��  �у�]� ������������̡hf�PH���  Q�Ѓ�������������U��hf�PH�EPQ���  �у�]� ̡hf�PH���   j Q�Ѓ�����������U��hf�PH�EPj Q���   �у�]� ��������������̡hf�PH���   jQ�Ѓ�����������U��hf�PH�EPjQ���   �у�]� ��������������̡hf�PH���   jQ�Ѓ����������U��hf�PH�EPjQ���   �у�]� ���������������U��hf�PH�EP�EPQ���   �у�]� �������������U��hf�PH�EP�EPQ���   �у�]� ������������̡hf�PH���   Q�Ѓ�������������U��hf�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���@���������t�E�hf�QH���   PVW�у���_^]� �����U��EVW���MPQ�L���������t�M�hf�BH���   QVW�҃���_^]� ̡hf�PH���   Q�Ѓ������������̡hf�PH���   Q�Ѓ�������������U��hf�PH�EPQ���   �у�]� �U��hf�PH�EPQ���   �у�]� �U��hf�PH�EP�EPQ��8  �у�]� �������������U��hf�PH�EP�EPQ��   �у�]� ������������̡hf�PH���  Q�Ѓ������������̡hf�PH���  Q�Ѓ������������̡hf�PH���  Q�Ѓ������������̡hf�PH��  Q�Ѓ������������̡hf�PH��  Q�Ѓ�������������U��hf�PH�EP�EPQ��  �у�]� �������������U��hf�PH�EP�EP�EPQ��   �у�]� ���������U��hf�PH�EP�EP�EP�EPQ��|  �у�]� �����U��hf�PH�EPQ��  �у�]� ̡hf�PH��T  Q�Ѓ�������������U��hf�PH�EP�EPQ��  �у�]� �������������U��hf�PH�EPQ��8  �у�]� �U��hf�PH�EPQ��<  �у�]� �U��hf�PH�EP�EP�EPQ��@  �у�]� ���������U��hf�PH�EPQ���  �у�]� ̡hf�PH��L  Q��Y��������������U��hf�PH�EPQ��H  �у�]� ̡hfV��H@�Q,WV�ҋhf�Q��j �ȋ��   h�  �Ћhf�QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡hf�P@�B,Q�Ћhf�Q��j �ȋ��   h�  �������U��hf�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��hf�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��hf�PH�EP�EP�EPQ��   �у�]� ��������̡hf�HH��  ��U��hf�HH��  ]��������������U��hf�E�PH��$  ���$Q�Ѓ�]� �����������̡hf�PH��(  Q�Ѓ�������������U��hf�PH�EP�EPQ��,  �у�]� �������������U��hf�E�PH�EP�E���$PQ��0  �у�]� ���̡hf�PH���  Q�Ѓ������������̡hf�PH��4  Q�Ѓ������������̋��     �������̡hf�PH���|  jP�у���������U��hf�UV��HH��x  R��3Ƀ������^��]� ��̡hf�PH���|  j P�у��������̡hf�PH��P  Q�Ѓ������������̡hf�PH��T  Q�Ѓ������������̡hf�PH��X  Q�Ѓ�������������U��hf�PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡hf�PH��`  Q�Ѓ�������������U��hf�PH�EPQ��d  �у�]� �U��hf�E�PH��h  ���$Q�Ѓ�]� ������������U��hf�E�PH��t  ���$Q�Ѓ�]� ������������U��hf�E�PH��l  ���$Q�Ѓ�]� ������������U��hf�PH�EPQ��p  �у�]� �U��hf�PH�EP�EP�EP�EPQ���  �у�]� �����U��hf�PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U��hf�E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E�hf�HH�E���   R�U���$P�ERP�у�]����������������U���E�M��$�|�  �M;�|�M;�~��]�����������U��hf�PH�E���   Q�MPQ�҃�]� ������������̡hf�PH���   Q��Y�������������̡hf�PH���   Q�Ѓ������������̡hf�PH���   Q��Y��������������U��hf�PH�EP�EPQ���   �у�]� �������������U��hf�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡hf�PH��t  Q��Y�������������̋�� �$�@    ���$�hf�Pl�A�JP��Y��������U��hfV��Hl�V�AR�ЋE����u
�   ^]� �hf�Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uËhf�QlP�B�Ѓ�������U��hf�Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E�hf�HH�ER�U���$P���  R�Ѓ�]����U��hf�HH���  ]��������������U��hf�HH���  ]��������������U��U0�E(�hf�HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U��hf�HH���  ]��������������U��hf�E�PH�EP���$Q���  �у�]� ��������U���SV����  �؉]����   �} ��   �hf�HH��p  j h�  V�҃��E��u
^��[��]� �MW3��}�� �  ����   �]��I �E�P�M�Q�MW还  ��ta�u�;u�Y�I ������u�E�������L�;Ht-�hf�Bl�S�@����QR�ЋD������t	�M�P裗  F;u�~��}��MG�}��n�  ;��v����]�_^��[��]� ^3�[��]� ��������������U����hfSV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u�hf�HH���  �'��u�hf�HH���  ���ušhf�HH���  S�ҋȃ��E��t�W�4�  �hf�HH���   h�  S3��҃����  ���_�u����    �hf�Hl�U�B�IWP�ы�������   �hf�F�J\�UP�A,R�Ѓ���t�K�Q�M�U�  �hf�F�J\�UP�A,R�Ѓ���t�K�Q�M�,�  �E��;Pt&�F�hf�Q\�J,P�EP�у���t	�MS���  �hf�v�B\�M�P,VQ�҃���t�M�CP�ӕ  �hf�QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U��hf�HH���   ]�������������̡hf�PH���   Q��Y��������������U��hf�HH���  ]��������������U��hf��P���   V�uW�}���$V�����E������At���E������z����؋hf�Q�B,���$V����_^]����������������U���0��hf�U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١hf�]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U��hf�HH�]��U��hf�H@�AV�u�R�Ѓ��    ^]�������������̡hf�HH�h�  �҃�������������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�HH�Vh  �ҋ�������   �EPh�  ��������t]�hf�QHj P���   V�ЋMQh(  �V�������t3�hf�JH���   j PV�ҡhf���   �B��j j���Ћ�^]áhf�H@�QV�҃�3�^]�������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�HH�Vh�  �ҋ�����u^]áhf�HH�U�E��  RPV�у���u�hf�B@�HV�у�3���^]�������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�HH�I]�����������������U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�PH�EPQ���  �у�]� �U��hf�PH�EPQ���  �у�]� ̡hf�PH���  Q�Ѓ�������������U��hf�HH���  ]��������������U��hf�E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡hf�PH���  Q�Ѓ�������������U��hf�PH�EP�EPQ���  �у�]� ������������̡hf�PH��  Q�Ѓ�������������U��hf�PH�EP�EP�EPQ���  �у�]� ��������̡hf�PH���  Q�Ѓ������������̡hf�PH���  Q�Ѓ�������������U��hf�PH�EPQ��  �у�]� �U��hf�PH�EPQ��  �у�]� ̋������������������������������̡hf�HH���  ��U��hf�HH���  ]��������������U��hf�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U��hf�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡hf�PH��,  Q�Ѓ�������������U��hf�PH�EPQ��X  �у�]� ̡hf�PH��\  Q�Ѓ�������������U��hf�HH��0  ]��������������U��hf��W���HH���   j h�  W�҃��} u�   _��]� Vh�  �������������   �hf�HH���   j VW�҃��M���L  �hf�P�E�R0Ph�  �M����E�hf�P�B,���$h�  �M��Ћhf�Q@�J(j �E�PV�у��M���L  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7�hf�U�HH���   RW�Ѓ���u�hf�QH���   jW�Ѓ���t�   �����   �hf�QH���   W�Ѓ��} u(�hf�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;�hf�U�HH�ER�USP���  VRW�Ћhf���   �B(�����Ћ���uŃ; u�hf�QH���   W�Ѓ���t3���   �W��u1�hf�QH���   �Ћhf�E�QH���   PW�у�_^[]� �hf�BH���   �у��} u0�hf�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� �hf�QH�h  �Ћ؃���u_^[]� �hf���   �u�Bx���Ћhf���   P�B|���Ѕ�tU�hf�E�QH�MP�Ej Q���  VPW�у���t�hf���   �ȋBHS�Ћhf���   �B(���Ћ���u�_^��[]� ��������������U��EV���u�hf�HH���  �'��u�hf�HH���  ���u�hf�HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D�hf�HH���   S�]VWh�  S�ҋ�hf�HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��.
  �hf���   �B���Ћhf=�  ��  �QH���   Wh:  S�Ћhf�QH�E����   h�  S�Ћhf�QHW�����   h�  S�uԉ}��Ћhf�QH�E苂  S�Ћhf�QH�EЋ��  S�Ѓ�(�E��E��$��~~�M���M�I �MЅ�tMj�W�A�  ���t@�@�Ẽ|� �4�~����%�������;�u/���p�  ;E�~�E؋��1�  E���E�;Pu�E���E��E�G;}�|��}� tv�u�j S�����������  ���������tV�������}�;�uK�hf�H���  �4�h�$��h�  V�҃��E���N  �M�PVP����P���  ����}ܡhf�H���  �4�h�$��h�  V�҃��E����  �M�3�;�t;�tVQP��  ���E�;�~-�hf�Qh�$��h�  P���   �Ѓ��E�;���  �hf�E��QH��  j�PS�у�����  �u�;�tjS����������{  ��������E���}�hf�BH���   Wh�  S�у�3�9}ԉE�}��`  �}���}Ȑ�MЅ��R  �U�j�R�J�  ����>  �M̍@�|� ���]�~����%�������9E���  ���=�  �E�3�3�9C�E܉M���   ��$    �����������tk�]��}������������ϋ9�<��}�@�҉��y�]��|��]�@@�z�<��y�]��|��]�@@�z�<��I�}��]�@���M��}�@����@�M�A;K�M��t����E؅��9  �+U�j��PR�M�赍  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$�$� �U����4�"�M����t��U����t�
�M����t�M���;]�|��E܃�F;]؉M��	����U�;U��
  �U�R��l  �E�P��l  �M�Q�l  ��_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���P�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@��;EԉE��}�������U�R�j  �E�P�j  ���  ���   �B����=  ��  �hf�QH���   j h(  S�Ћhf�QH�����   h(  S�ЋЃ�3��U؅�~'����    �ǅ�t�|� t�4N��tN�@;�|�u��u܋hf�Q���  �4v�h�$��hK  V�Ѓ��E�����   �M��t��tVQP��  ���u؋hf�Q���  �h�$��hP  V�Ѓ��E���tP��t��tVWP�ֳ  ���M����+hf�RH��PQ�E���   S�Ѓ���u�M�Q�bi  �U�R�Yi  ��_^3�[��]áhf�HH���   j h�  S�҉E��hf�HH���   j h(  S��3�3���3�9]؉E��}ĉ]��7  �U��څ��  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�F@F����;�|��}ă|� ts�U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�F�v�Ћ��A�B�A�B�A�B�A�B�I�J�U�F<ډ}�C;]؉]�������M�3�3�;�~�U����$    ��t���   @;�|��U�R�g  ���E�P�g  ��_^�   [��]�o� z� �� �� ������������U��E� �M+]� ���������������U��V��V��$�hf�Hl�AR�Ѓ��Et	V�Tj  ����^]� ����������U��hf�P8�EPQ�JD�у�]� ���̡hf�H8�Q<�����U��hf�H8�A@V�u�R�Ѓ��    ^]�������������̡hf�H8�������U��hf�H8�AV�u�R�Ѓ��    ^]��������������U��hf�P8�EP�EP�EPQ�J�у�]� ������������U��hf�P8�EP�EPQ�J�у�]� �hf�P8�BQ�Ѓ����������������U��hf�P8�EPQ�J �у�]� ����U��hf�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U��hf�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U��hf�P8�EP�EPQ�J(�у�]� U��hf�P8�EP�EP�EPQ�J,�у�]� ������������U��hf�P8�EP�EP�EPQ�J�у�]� ������������U��hf�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U��hf�P8�EP�EPQ�J0�у�]� U��hf�P8�EP�EP�EPQ�J4�у�]� ������������U��hf�P8�EPQ�J8�у�]� ����U��hf�H��x  ]��������������U��hf�H��|  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H�A,]�����������������U��hf�H���  ]��������������U��hf�H�QV�uV�ҡhf�H�Q8V�҃���^]�����̡hf�H�Q<�����U��hf�H�I@]����������������̡hf�H�QD����̡hf�H�QH�����U��hf�H�AL]�����������������U��hf�H�IP]�����������������U��hf�H��<  ]��������������U��hf�H��,  ]��������������U��hf�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡hf�H���   ��hf�H���  ��U��hf�H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U��hf�H�A]�����������������U��hf�H��\  ]��������������U��hf�H�AT]�����������������U��hf�H�AX]�����������������U��hf�H�A\]����������������̡hf�H�Q`�����U��hf�H���  ]�������������̡hf�H�Qd����̡hf�H�Qh�����U��hf�H�Al]�����������������U��hf�H�Ap]�����������������U��hf�H�At]�����������������U��hf�H��D  ]��������������U��hf�H��  ]��������������U��hf�H�Ix]�����������������U��hf�H��@  ]��������������U��V�u���B  �hf�H�U�A|VR�Ѓ���^]���������U��hf�H���   ]��������������U��hf�H��h  ]��������������U��hf�H��d  ]��������������U��hf�H���  ]�������������̡hf�H���   ��U��hf�H��l  ]��������������U��hf�H��   ]��������������U��hf�H��  ]��������������U��V�u���6  �hf�H���   V�҃���^]���������̡hf�H��`  ��U��hf�H��  ]��������������U��hf�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U��hf�H���  ]��������������U��U�E�hf�H�E���   R���\$�E�$P�у�]�U��hf�H���   ]��������������U��hf�H���   ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���   ]��������������U��hf�H���   ]��������������U��hf�H���   ]��������������U��hf�H���   ]��������������U��hf�H���   ]��������������U��hf�H���   ]��������������U��hf�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��hf�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��hf�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��hf�H��8  ]��������������U��V�u(V�u$�E�@�hf�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@�hf�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��hf�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U��hf�P0�EP�EP�EP�EPQ���   �у�]� ����̡hf�P0���   Q�Ѓ�������������U��hf�P0�EP�EPQ���   �у�]� �������������U��hf�P0�EP�EP�EP�EPQ���   �у�]� ����̡hf�P0���   Q�Ѓ������������̡hf�H0���   ��U��hf�H0���   V�u�R�Ѓ��    ^]�����������U��hf�H��H  ]��������������U��hf�H��T  ]�������������̡hf�H��p  ��hf�H���  ��U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �hf���   �Qj PV�ҡhf���   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M��
0  P�E�hicMCP�k������M��00  �hf���   �JT�E�P�у���u(�u���/  �hf���   ��M�Q�҃���^��]áhf���   �AT�U�R�Ћu��P���/  �hf���   �
�E�P�у���^��]�������������U��hf�H��  ]��������������U��hf�H��\  ]��������������U��hf�H�U��t  ��V�uVR�E�P�у����  �M��K  ��^��]�����U��hf�H�U���  ��VWR�E�P�ыhf�u���B�HV�ыhf�B�HVW�ыhf�B�P�M�Q�҃�_��^��]����������������U��hf�H�U���  ��VWR�E�P�ыhf�u���B�HV�ыhf�B�HVW�ыhf�B�P�M�Q�҃�_��^��]����������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H�U�E��VWj R�UP�ERP��t  �U�R�Ћhf�Q�u���BV�Ћhf�Q�BVW�Ћhf�Q�J�E�P�у�(_��^��]��U��hf�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �hf���   j P�BV�Ћhf���   �
�E�P�у�$��^��]���U��hf�H��8  ]��������������U���  � Q3ŉE��M�EPQ������h   R��  ����|	=�  |#��hf�H��0  h�$hH  �҃��E� �hf�H��4  ������Rh,%�ЋM�3̓����  ��]�������U��hf�H��  ��V�U�WR�Ћhf�Q�u���BV�Ћhf�Q�BVW�Ћhf�Q�J�E�P�у�_��^��]����U��hf�H��  ��V�U�WR�Ћhf�Q�u���BV�Ћhf�Q�BVW�Ћhf�Q�J�E�P�у�_��^��]����U��hf�H��p  ��$�҅�trh���M���*  �hf�P�E�R4Ph���M��ҡhf�P�E�R4Ph���M���j �E�P�M�hicMCQ�����hf���   ��M�Q�҃��M���*  ��]�U��hf�H��p  ��$V�҅�u�hf�H�u�QV�҃���^��]�Wh!���M��<*  �hf�P�E�R4Ph!���M���j �E�P�M�hicMCQ�����hf���   �QHP�ҋu���hf�H�QV�ҡhf�H�QVW�ҡhf���   ��U�R�Ѓ�$�M���)  _��^��]������U��hf�H��p  ��$V�҅�u�hf�H�u�QV�҃���^��]�Wh����M��l)  �hf�P�E�R4Ph����M���j �E�P�M�hicMCQ�����hf���   �QHP�ҋu���hf�H�QV�ҡhf�H�QVW�ҡhf���   ��U�R�Ѓ�$�M��-)  _��^��]������U��hf�H��p  ��$�҅�u��]�Vh#���M��(  �hf�P�E�R4Ph#���M���j �E�P�M�hicMCQ������hf���   �Q8P�ҋ�hf���   ��U�R�Ѓ��M��(  ��^��]���������������U��hf�H��p  ��$�҅�u��]�Vhs���M��(  �hf�P�E�R4Phs���M���j �E�P�M�hicMCQ�W����hf���   �Q8P�ҋ�hf���   ��U�R�Ѓ��M���'  ��^��]���������������U��hf�H���  ]��������������U��hf�H��@  ]��������������U��hf�H���  ]��������������U��V�u���t�hf�QP��D  �Ѓ��    ^]������U��hf�H��H  ]��������������U��hf�H��L  ]��������������U��hf�H��P  ]��������������U��hf�H��T  ]��������������U��hf�H��X  ]��������������U��hf�H��\  ]�������������̡hf�H��d  ��U��hf�H��h  ]��������������U��hf�H��l  ]�������������̡hf�H���  ��U��hf�H�U���  ��VR�E�P�ыu��P����%  �M���%  ��^��]�����U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H��l  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H��$  ]��������������U��hf�H��(  ]��������������U��hf�H��,  ]�������������̡hf�H��0  ��hf�H��<  ��U��hf�H���  ]�������������̡hf�H���  ��U��hf�H���  ]������������������������������U��hf�H��  ]�������������̡hf�H��P  ��U��hf�H��`  ]�������������̡hf���   ���   ��Q��Y��������U��hf�H�A�U��� R�Ћhf�Q�Jj j��E�h0%P�ыUR�E�P�M�Q�����hf�B�P�M�Q�ҡhf�H�A�U�R�Ћhf�Q�J�E�P�у�,��]��U��hf�P�EP�EP�EPQ�J�у�]� �����������̡hfV��H�QV�ҡhf�H$�QDV�҃���^�����������U��hfV��H�QV�ҡhf�H$�QDV�ҡhf�U�H$�AdRV�Ѓ���^]� ��U��hfV��H�QV�ҡhf�H$�QDV�ҡhf�U�H$�ARV�Ѓ���^]� ��U��hfV��H�QV�ҡhf�H$�QDV�ҡhf�H$�U�ALVR�Ѓ���^]� �̡hfV��H$�QHV�ҡhf�H�QV�҃�^�������������U��hf�P$�EPQ�JL�у�]� ����U��hf�P$�R]�����������������U��hf�P$�Rl]����������������̡hf�P$�Bp����̡hf�P$�BQ�Ѓ����������������U��hf�P$��VWQ�J�E�P�ыhf�u���B�HV�ыhf�B�HVW�ыhf�B�P�M�Q�҃�_��^��]� ���U��hf�P$�EPQ�J�у�]� ����U��hf�P$��VWQ�J �E�P�ыhf�u���B�HV�ыhf�B$�HDV�ыhf�B$�HLVW�ыhf�B$�PH�M�Q�ҡhf�H�A�U�R�Ѓ� _��^��]� ���U��hf�P$��VWQ�J$�E�P�ыhf�u���B�HV�ыhf�B$�HDV�ыhf�B$�HLVW�ыhf�B$�PH�M�Q�ҡhf�H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e����hf�Q$�JH�E�P�ыhf�B�P�M�Q�҃���^��]� ����̡hf�P$�B(Q��Yáhf�P$�BhQ��Y�U��hf�P$�EPQ�J,�у�]� ����U��hf�P$�EPQ�J0�у�]� ����U��hf�P$�EPQ�J4�у�]� ����U��hf�P$�EPQ�J8�у�]� ����U��hf�UV��H$�ALVR�Ѓ���^]� ��������������U��hf�H�QV�uV�ҡhf�H$�QDV�ҡhf�H$�U�ALVR�Ћhf�E�Q$�J@PV�у���^]�U��hf�UV��H$�A@RV�Ѓ���^]� ��������������U��hf�P$�EPQ�J<�у�]� ����U��hf�P$�EPQ�J<�у����@]� ���������������U��hf�P$�EP�EPQ�JP�у�]� U��hf�P$�EPQ�JT�у�]� ���̡hf�H$�QX�����U��hf�H$�A\]�����������������U��hf�P$�EP�EP�EPQ�J`�у�]� �����������̡hf�H(�������U��hf�H(�AV�u�R�Ѓ��    ^]��������������U��hf�P(�R]����������������̡hf�P(�B�����U��hf�P(�R]�����������������U��hf�P(�R]�����������������U��hf�P(�R ]�����������������U��hf�P(�E�RjP�EP��]� ��U��hf�P(�E�R$P�EP�EP��]� �hf�P(�B(����̡hf�P(�B,����̡hf�P(�B0�����U��hf�P(�R4]�����������������U��hf�P(�RX]�����������������U��hf�P(�R\]�����������������U��hf�P(�R`]�����������������U��hf�P(�Rd]�����������������U��hf�P(�Rh]�����������������U��hf�P(�Rl]�����������������U��hf�P(�Rx]�����������������U��hf�P(���   ]��������������U��hf�P(�Rt]�����������������U��hf�P(�Rp]�����������������U��hf�P(�BpVW�}W���Ѕ�t:�hf�Q(�Rp�GP���҅�t"�hf�P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U��hf�P(�BtVW�}W���Ѕ�t:�hf�Q(�Rt�GP���҅�t"�hf�P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U��VW�}W���0�����t8�GP���!�����t)�OQ��������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W���0�����t8�GP���!�����t)�O0Q��������t��HW��������t_�   ^]� _3�^]� ������������U����hf�E�    �E�    �P(�RhV�E�P���҅���   �E���uG�hf�H�A�U�R�Ћhf�Q�E�RP�M�Q�ҡhf�H�A�U�R�Ѓ��   ^��]� �hf�Qh4%he  P���   �Ћhf���E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P��?  ��3�^��]� �M��U�j IQ�MR������E�P��?  ���   ^��]� ���������������U��hf��V��H�A�U�R�Ѓ��M�Q������^��u�hf�B�P�M�Q�҃�3���]� �hf�H$�E�I�U�RP�ыhf�B�P�M�Q�҃��   ��]� �U��Q�hf�P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U��hf�P(�R8]�����������������U��hf�P(�R<]�����������������U��hf�P(�R@]�����������������U��hf�P(�RD]�����������������U��hf�P(�RH]�����������������U��hf�P(�E�R|P�EP��]� ����U��hf�P(�RL]�����������������U��hf�E�P(�BT���$��]� ���U��hf�E�P(�BPQ�$��]� ����̡hf�H(�Q�����U��hf�H(�AV�u�R�Ѓ��    ^]��������������U��hf�P(���   ]��������������U��hf�H(�A]����������������̡hf�H,�Q,����̡hf�P,�B4�����U��hf�H,�A0V�u�R�Ѓ��    ^]�������������̡hf�P,�B8�����U��hf�P,�R<��VW�E�P�ҋu���hf�H�QV�ҡhf�H$�QDV�ҡhf�H$�QLVW�ҡhf�H$�AH�U�R�Ћhf�Q�J�E�P�у�_��^��]� �������U��hf�P,�E�R@��VWP�E�P�ҋu���hf�H�QV�ҡhf�H�QVW�ҡhf�H�A�U�R�Ѓ�_��^��]� ��̡hf�H,�j j �҃��������������U��hf�P,�EP�EPQ�J�у�]� U��hf�H,�AV�u�R�Ѓ��    ^]�������������̡hf�P,�B����̡hf�P,�B����̡hf�P,�B����̡hf�P,�B ����̡hf�P,�B$����̡hf�P,�B(�����U��hf�P,�R]�����������������U��hf�P,�R��VW�E�P�ҋu���hf�H�QV�ҡhf�H$�QDV�ҡhf�H$�QLVW�ҡhf�H$�AH�U�R�Ћhf�Q�J�E�P�у�_��^��]� �������U��hf�H��D  ]��������������U��hf�H��H  ]��������������U��hf�H��L  ]��������������U��hf�H�I]�����������������U��hf�H�A]�����������������U��hf�H�I]�����������������U��hf�H�A]�����������������U��hf�H�I]�����������������U��hf�H���  ]��������������U��hf�H�A]�����������������U���V�u�E�P��������hf�Q$�J�E�P�у���u-�hf�B$�PH�M�Q�ҡhf�H�A�U�R�Ѓ�3�^��]Ëhf�Q�J�E�jP�у���u=�U�R��������u-�hf�H$�AH�U�R�Ћhf�Q�J�E�P�у�3�^��]Ëhf�B�HjV�у���u�hf�B�HV�у����I����hf�Q$�JH�E�P�ыhf�B�P�M�Q�҃��   ^��]�����������U��hf�H�A ]�����������������U��hf�H�I(]�����������������U��hf�H��  ]��������������U��hf�H��   ]��������������U��hf�H��  ]��������������U��hf�H��  ]��������������U��hf�H�A$��V�U�WR�Ћhf�Q�u���BV�Ћhf�Q$�BDV�Ћhf�Q$�BLVW�Ћhf�Q$�JH�E�P�ыhf�B�P�M�Q�҃�_��^��]������U��hf�H���  ��V�U�WR�Ћhf�Q�u���BV�Ћhf�Q$�BDV�Ћhf�Q$�BLVW�Ћhf�Q$�JH�E�P�ыhf�B�P�M�Q�҃�_��^��]���U��hf�H���  ]��������������U���<��fSVW�E�    ��t�E�P�   �������/�hf�Q�J�E�P�   �ыhf�B$�PD�M�Q�҃��}�hf�H�u�QV�ҡhf�H$�QDV�ҡhf�H$�QLVW�҃���t)�hf�H$�AH�U�R����Ћhf�Q�J�E�P�у���t&�hf�B$�PH�M�Q�ҡhf�H�A�U�R�Ѓ�_��^[��]���U��hf�H�U���  ��VWR�E�P�ыhf�u���B�HV�ыhf�B$�HDV�ыhf�B$�HLVW�ыhf�B$�PH�M�Q�ҡhf�H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]����������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]��������������U��hf�H���  ]�������������̡hf�H���   ��U��hf�H���   V�uV�҃��    ^]�������������U��hf�P�]��hf�P�B����̡hf�P���   ��U��hf�P�R`]�����������������U��hf�P�Rd]�����������������U��hf�P�Rh]�����������������U��hf�P�Rl]�����������������U��hf�P�Rp]�����������������U��hf�P�Rt]�����������������U��hf�P���   ]��������������U��hf�P��  ]��������������U��hf�P�Rx]�����������������U��hf�P���   ]��������������U��hf�P�R|]�����������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P�EPQ��  �у�]� �U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��E��t �hf�R P�B$Q�Ѓ���t	�   ]� 3�]� U��hf�P �E�RLQ�MPQ�҃�]� U��E��u]� �hf�R P�B(Q�Ѓ��   ]� ������U��hf�P�R]�����������������U��hf�P�R]�����������������U��hf�P�R]�����������������U��hf�P�R]�����������������U��hf�P�R]�����������������U��hf�P�R]�����������������U��hf�P�E�R\P�EP��]� ����U��hf�P�E��  P�EP��]� �U��hf�E�P�B ���$��]� ���U��hf�E�P�B$Q�$��]� �����U��hf�E�P�B(���$��]� ���U��hf�P�R,]�����������������U��hf�P�R0]�����������������U��hf�P�R4]�����������������U��hf�P�R8]�����������������U��hf�P�R<]�����������������U��hf�P�R@]�����������������U��hf�P�RD]�����������������U��hf�P�RH]�����������������U��hf�P�RL]�����������������U��hf�P�RP]�����������������U��hf�P���   ]��������������U��hf�P�RT]�����������������U��hf�P�EPQ��  �у�]� �U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P�RX]����������������̡hf�P���   ��U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]��������������U��hf�P���   ]�������������̡hf�P���   ��U��hf�P���   ]�������������̡hf�P���   ��hf�P���   ��hf�P���   ��U��hf�H���   ]��������������U��hf�H��   ]��������������U��hf�H�U�E��VWRP���  �U�R�Ћhf�Q�u���BV�Ћhf�Q�BVW�Ћhf�Q�J�E�P�у�_��^��]������������U��hf�H���  ]��������������U��hf�P(�BPVW�}�Q�]���E�$�Ѕ�tM�hf�G�Q(�]�E�BPQ���$�Ѕ�t,�hf�G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U��hf�P(�BTVW�}����$���Ѕ�tE�hf�G�Q(�BT�����$�Ѕ�t(�hf�G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U��hf�P(�} �R8����P��]� �U��hf�P�BdS�]VW��j ���Ћhf�Q�����   h4%Fh�  V�Ћhf���E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћhf�Q(�BHV���Ѕ�t �hf�Q(�E�R VP���҅�t�   �3��EP�(  ��_��^[]� ������U���V�E���MP�k���P���#����hf�Q�J���E�P�у���^��]� ��̡hf�P�BVj j����Ћ�^���������U��hf�P�E�RVj P���ҋ�^]� U��hf�P�E�RVPj����ҋ�^]� �hf�P�B�����U��hf�P���   Vj ��Mj V�Ћ�^]� �����������U��hf�P�EPQ�J�у�]� ����U��hf�P�EPQ�J�у����@]� ���������������U��hf�P�E�RtP�ҋhf���   P�BX�Ѓ�]� ���U��hf�P�E�Rlh#  P�EP��]� ���������������U��hf�P�E�RlhF  P�EP��]� ���������������U��hf�P�E�RtP�ҋhf���   �M�R`QP�҃�]� ���������������U��hf�P���   ]��������������U��hf�P�E���   P�҅�u]� �hf���   P�B�Ѓ�]� �������̡hf�HL���   ��U��hf�H@�AV�u�R�Ѓ��    ^]�������������̡hf�HL�������U��hf�H@�AV�u�R�Ѓ��    ^]�������������̡hf�PL���   Q�Ѓ�������������U��hf�PL�EP�EPQ���   �у�]� �������������U��hfV��HL���   V�҃���u�hf�U�HL���   j RV�Ѓ�^]� �hf���   �ȋBP�Ћhf���   �MP�BH��^]� �����̡hf�PL��(  Q�Ѓ�������������U��hf�PL�EP�EPQ��,  �у�]� ������������̡hf�HL�Q�����U��hf�H@�AV�u�R�Ѓ��    ^]��������������U��hf�PL�E�R��VPQ�M�Q�ҋu��P���%����M��=�����^��]� ����U��hf�PL�EPQ���   �у�]� �U��hf�PL�EP�EPQ�J�у�]� �hf�PL�BQ�Ѓ���������������̡hf�PL�BQ�Ѓ���������������̡hf�PL�BQ�Ѓ����������������U��hf�PL�EP�EP�EPQ�J �у�]� ������������U��hf�PL�EPQ��4  �у�]� �U��hf�PL�EP�EP�EPQ�J$�у�]� ������������U��hf�PL�EP�EP�EP�EPQ�J(�у�]� �������̡hf�PL�B,Q�Ѓ���������������̡hf�PL�B0Q�Ѓ����������������U��hf�PL�EP�EPQ��  �у�]� ������������̡hf�PL���   Q�Ѓ�������������U��hf�PL�E��  ��VPQ�M�Q�ҋu��P�������M�������^��]� ̡hf�PL�B4Q�Ѓ���������������̡hf�PL�B8j Q�Ѓ��������������U��hf�PL���   ]��������������U��hf�PL���   ]��������������U��hf�PL���   ]��������������U��hf�PL���   ]��������������U��hf�PL���   ]��������������U��hf�PL���   ]��������������U��hf�PL��l  ]��������������U��hf�PL���   ]��������������U��hf�PL���   ]��������������U��hf�PL���   ]��������������U��hf�PL�EPQ�J<�у�]� ���̡hf�PL�BQ��Y�U��hf�PL�EP�EPQ�J@�у�]� U��hf�PL�Ej PQ�JD�у�]� ��U��hf�PL�Ej PQ�JH�у�]� ��U��hf�PL�EjPQ�JD�у�]� ��U��hf�PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��4{��W�M�Q�U�R���������M����'m����t�hf���   ��U�R�Ѓ�_^3�[��]Ëhf���   �J8�E�P�ыhf�����   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  �~z��j�M�Q�U�R���]����M��ul���hf���   ��U�R�Ѓ�^��]�����������U���$�hf�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}���y��j�E�P�M�Q���ف���M���k���hf���   ��M�Q�҃�_^��]� ��U���$�hf�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��zy��j�E�P�M�Q���Y����M��qk���hf���   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��y��W�M�Q�U�R���Ԁ�����M����k����t+�u���y����hf���   ��U�R�Ѓ�_��^[��]� �hf���   �JL�E�P�ыu��P��������hf���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��Tx��W�M�Q�U�R���������M����Gj����t+�u�������hf���   ��U�R�Ѓ�_��^[��]� �hf���   �JL�E�P�ыu��P���%����hf���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��w��W�M�Q�U�R���T�����M����i��_^��[t�hf���   ��U�R�������]Ëhf���   �J<�E�P���]��hf���   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}���v��W�M�Q�U�R���~�����M�����h����t�hf���   ��U�R�Ѓ�_^3�[��]Ëhf���   �J8�E�P�ыhf�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��4v��W�M�Q�U�R����}�����M����'h����t-��u�hf����   ���^�U�R�Ѓ�_��^[��]� �hf���   �JP�E�P�ы�u�H��P�@�N�hf�V���   �
�F�E�P�у�_��^[��]� �����̡hf�PL���   Q��Y��������������U��hf�PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U��hf�PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��t��W�M�Q�U�R���d|�����M����f����t-��u�hf����   ���^�U�R�Ѓ�_��^[��]� �hf���   �JP�E�P�ы�u�H��P�@�N�hf�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���s��W�M�Q�U�R���{�����M�����e����t-��u�hf����   ���^�U�R�Ѓ�_��^[��]� �hf���   �JP�E�P�ы�u�H��P�@�N�hf�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��s��W�M�Q�U�R����z�����M�����d����t-��u�hf����   ���^�U�R�Ѓ�_��^[��]� �hf���   �JP�E�P�ы�u�H��P�@�N�hf�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��4r��W�M�Q�U�R����y�����M����'d����t�hf���   ��U�R�Ѓ�_^3�[��]Ëhf���   �J8�E�P�ыhf�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  �q��j�M�Q�UR���^y���M�vc���hf���   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��q��j�U�R�E�P����x���M��c���hf���   �
�E�P�у�^��]� ��������U���$�hf�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��p��j�E�P�M�Q���ix���M��b���hf���   ��M�Q�҃�_^��]� ��U���$�hf�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
p��j�E�P�M�Q����w���M��b���hf���   ��M�Q�҃�_^��]� ��U���$�hf�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��o��j�E�P�M�Q���iw���M��a���hf���   ��M�Q�҃�_^��]� ��U���$�hf�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
o��j�E�P�M�Q����v���M��a���hf���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��n��j�U�R�E�P���~v���M��`���hf���   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}��4n��W�M�Q�U�R����u�����M����'`����t-��u�hf����   ���^�U�R�Ѓ�_��^[��]� �hf���   �JP�E�P�ы�u�H��P�@�N�hf�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��dm��W�M�Q�U�R���$u�����M����W_����t�hf���   ��U�R�Ѓ�_^3�[��]Ëhf���   �J8�E�P�ыhf�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��l��W�M�Q�U�R���tt�����M����^����t�hf���   ��U�R�Ѓ�_^3�[��]Ëhf���   �J8�E�P�ыhf�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ���̡hf�PL���  ��U���$�hf�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��k��j�E�P�M�Q���s���M��]���hf���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��Ok��j�U�R�E�P���.s���M��F]���hf���   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���j��j�U�R�E�P���r���M���\���hf���   �
�E�P�у�^��]� ��������U��hf�H���   ]��������������U��hf�H���   ]�������������̡hf�H���   ��hf�H���   ��U��hf�H���   V�u�R�Ѓ��    ^]�����������U��hf�H���   ]��������������U��hf�HL�QV�ҋ���u^]áhf�H�U�Ej R�UP��h  RV�Ѓ���u�hf�Q@�BV�Ѓ�3���^]��������U��hf�H�U�E��h  j R�U�� P�ERP�у�]����U��hf�H���   ]��������������U��hf�H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡hf�PL�BLQ�Ѓ���������������̡hf�PL�BPQ�Ѓ����������������U��hf�PL�EP�EPQ�JT�у�]� U��hf�PL�EPQ��  �у�]� �U��hf�PL�EPQ���   �у�]� ̡hf�PL�BXQ�Ѓ����������������U��hf�PL�EP�EP�EPQ�J\�у�]� ������������U���4�hfSV��HL�QW�ҋ�3ۉ}�;��x  �M�������hf�E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡhf���   �BSSW���Ѕ���   �hf�QL�BW�Ћ���;���   ��    �hf���   �B(���ЍM�Qh�   ���u��j���������   �M�;���   �hf���   ���   S��;�tm�hf���   �ȋB<V�Ћhf���   ���   �E�P�у�;�t�hf�B@�HV�у���;��\����}��M�聿���M�������_^[��]� �}��hf�B@�HW�ыhf���   ���   �M�Q�҃��M��9����M������_^3�[��]� �����̡hf�PL�B`Q�Ѓ���������������̡hf�PL�BdQ�Ѓ����������������U��hf�PL�EPQ�Jh�у�]� ���̡hf�PL��D  Q�Ѓ������������̡hf�PL�BlQ�Ѓ����������������U��hf�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh� h�� h�� h�� R�Q�U R�UR�UR�U���A�$�5hf�vLRP���   Q�Ѓ�4^]�  ������̡hf�PL���   Q�Ѓ�������������U��hf�PL�EP�EP�EPQ��   �у�]� ���������U��hf�PL��H  ]�������������̡hf�PL��L  ��U��hf�PL��P  ]��������������U��hf�PL��T  ]��������������U��hf�PL��p  ]��������������U��hf�PL��t  ]��������������U��hf�PL�EP�EP�EP�EP�EPQ���   �у�]� �U��hf�PL�EP�EP�EPQ���   �у�]� ���������U��hf�PL�EP�EP�EP�EPQ��   �у�]� �����U��hf�HL���   ]��������������U��hf�HL���   ]��������������U��hf�HL���   ]�������������̡hf�HL��  ��hf�HL��@  ��U��hf�PL���  ]��������������U��hf�PL���  ]��������������U��hf�PL���  ]��������������U��� �hfV3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\�hf�QLjP���   ���ЋM��U�Rh=���M�}��������hf���   ���   �U�R�Ѓ��M��u�茺����_^��]Ëhf���   ���   �E�P�у��M��u��^���_�   ^��]����U��� �hfV3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\�hf�QLjP���   ���ЋM��U�Rh<���M�}��C������hf���   ���   �U�R�Ѓ��M��u�輹����_^��]Ëhf���   ���   �E�P�у��M��u�莹��_�   ^��]����U���EV���V��������Au�hf�H��0  hx%j,�����^��^]� �����U���W������G���U���$������A�  ������A��   ��%������AuR������AuKV����M  ����M  �ȅ�u��^����__��]Ëƙ����ʅ�u�u��E�^������__��]���������Au������=�%��������Au6�����������U������G�����_��������Au�����U����_�
����������}Q  �E����U���%��������A{���������__��]�������������__��]����U����%V�E��������At����%������Au�������!����%�$�*Q  �����!���^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3�����%;���W���$���P  ��E����%�$�P  �V����������Au�hf�H��0  hx%j�����^����_u������������^]� ���U������EV�ы�������z!�hf�؋H��0  hx%j5�����U������$�	P  �]��F�$��O  �}��$��O  ��E�$��O  �^�����&���^��]� ��������������̋�� �%����������%���������̅�t��j�����̡hf�P��  ��hf�P��(  ��U��hf�P��   ��V�E�P�ҋuP���Z����M�蒷����^��]� ��������̡hf�P��$  ��U��hf�H��  ]��������������U��hf�H���  ]�������������̡hf�H��  ��U��hf�H���  ]��������������U��hf�H��x  ]��������������U��hf�H��|  ]�������������̡hf�H��d  ��U��hf�H��p  ]��������������U��hf�H��t  ]��������������U���EV����%t	V�X  ����^]� ��������������U��V�u���t�hf�QP��Ѓ��    ^]���������̡hf�H��@  hﾭ���Y����������U��E��t�hf�QP��@  �Ѓ�]����������������U��hf�H���  ]��������������U��hf�H��  ]�������������̡hf�H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�XN  ������u_^]Ã} tWj V�O  ��_������F�|f   ^]���U��hf�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW��M  ������u_^]�Wj V�N  ��_������F�|f   ^]�������������U��hf�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�\M  ������u_^]�Wj V�N  ��_������F�|f   ^]�������������U��hf�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW��L  ������u_^]�Wj V�M  ��_������F�|f   ^]�������������U��hf�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�\L  ������u_^]�Wj V�M  ��_������F�|f   ^]�������������U��M��t-�=|f t�y���A�uP�HM  ��]áhf�P�Q�Ѓ�]��������U��M��t-�=|f t�y���A�uP�M  ��]áhf�P�Q�Ѓ�]��������U��hf�H�U�R�Ѓ�]���������U��hf�H�U�R�Ѓ�]���������U��hf�E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�K  ������u_^]�Wj V��K  ��_������F�|f   ^]���������U��hf�E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   �hf��t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�)J  ������u_^]�Wj V��J  ��_������F�|f   ^]����������U��E��w�   �hf��t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�I  ������u_^]�Wj V�PJ  ��_������F�|f   ^]�������U��hf�H�U�R�Ѓ�]���������U��hf�H�U�R�Ѓ�]���������U��hf�H�U�R�Ѓ�]���������U��hf�H�U�R�Ѓ�]���������U��hf�P�E���   ��VWP�EP�E�P�ҋu���hf�H�QV�ҡhf�H�QVW�ҡhf�H�A�U�R�Ѓ�_��^��]� ������������U��E��u��f�MP�EPQ�cF����]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h�%j;h�fj��������t
W��螮���3��F��u_^]� �~ t3�9_��^]� �hf�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   �hf�H<�Q��3Ʌ����^��������������̃y t�   ËA��uËhf�R<P��JP�у��������U����u�hf�H�]� �hf�J<�URP�A�Ѓ�]� ���������������U�졀f��u�hf�H�]Ëhf�J<�URP�A�Ѓ�]�U�졀f��$V��u�hf�H�1��hf�J<�URP�A�Ѓ����hf�Q�J�E�SP�ыhf�B�P�M�QV�ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@�� j �M�Q�U�R�M��Ћhf�Q�J���E�P���у���[t.�hf�B�u�HV�ыhf�B�P�M�Q�҃���^��]áhf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M��ҡhf�H�u�QV�ҡhf�H�A�U�VR�Ћhf�Q�J�E�P�у���^��]���������������U�졀f��$SV��u�hf�H�1��hf�J<�URP�A�Ѓ����hf�Q�J�E�P�ыhf�B�P�M�QV�ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@�� j �M�Q�U�R�M��Ћhf�Q�J���E�P���у���t/�hf�B�u�HV�ыhf�B�P�M�Q�҃���^[��]áhf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M��ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@��j �M�Q�U�R�M��Ћhf�Q�J���E�P���у����3����hf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M��ҡhf�H�u�QV�ҡhf�H�A�U�VR�Ћhf�Q�J�E�P�у���^[��]����������������U�졀f��$SV��u�hf�H�1��hf�J<�URP�A�Ѓ����hf�Q�J�E�P�ыhf�B�P�M�QV�ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@�� j �M�Q�U�R�M��Ћhf�Q�J���E�P���у���t/�hf�B�u�HV�ыhf�B�P�M�Q�҃���^[��]áhf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M��ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@��j �M�Q�U�R�M��Ћhf�Q�J���E�P���у����3����hf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M��ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@��j �M�Q�U�R�M��Ћhf�Q�J���E�P���у���������hf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M��ҋu�E�P������hf�Q�J�E�P�у���^[��]�������U�졀f��$SV��u�hf�H�1��hf�J<�URP�A�Ѓ����hf�Q�J�E�P�ыhf�B�P�M�QV�ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@�� j �M�Q�U�R�M��Ћhf�Q�J���E�P���у���t/�hf�B�u�HV�ыhf�B�P�M�Q�҃���^[��]áhf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M��ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@��j �M�Q�U�R�M��Ћhf�Q�J���E�P���у����3����hf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M��ҡhf�H�A�U�R�Ћhf�Q�Jj j��E�h4&P�ыhf�B�@@��j �M�Q�U�R�M��Ћhf�Q�J���E�P���у���������hf�P�E��RHjP�M��ҡhf�P�E�M��RLj�j�PQ�M���j h4&�M��"���hf�P�R@j �E�P�M�Q�M��҅��hf�H�A�U�R���Ѓ���t/�hf�Q�u�BV�Ћhf�Q�J�E�P�у���^[��]Ëhf�M��B�PHjQ�M��ҡhf�P�E�M��RLj�j�PQ�M��ҋu�E�P���K���hf�Q�J�E�P�у���^[��]���������������U��hf�H<�A]����������������̡hf�H<�Q�����V��~ u>���t�hf�Q<P�B�Ѓ��    W�~��t���
���W�������F    _^��������U���V�E�P���>�����P��������M���ɣ����^��]��̃=�f uK��f��t�hf�Q<P�B�Ѓ���f    ��f��tV��耣��V�z�������f    ^������������U���8�hf�H�AS�U�V3�R�]��Ћhf�Q�JSj��E�h8&P�ыhf�B<�P�M�Q�ҋ�hf�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��2  �M�Q�U�R�M���2  ����   W�}�}���   �hf���   �U��ATR�Ћ�����tB�hf�Q�J�E�P���у��U�Rj�E�P�������hf�Q�ȋBxW���E���t�E� ��t�hf�Q�J�E�P����у���t�hf�B�P�M�Q����҃��}� u"�E�P�M�Q�M��2  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3ۉ]�;�u_�hf�H�A�U�R�Ћhf�Q�JSj��E�h8&P�ыhf�B<�P�M�Q�ҋ�hf�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��1  �M�Q�U�R�M��Q1  ���p  W�}��I �E����   �hf���   �U��ATR�Ћ�������   �hf�Q�J�E�P���ыhf�B���   ���M�Qj�U�R���Ћhf�Q�J���E�P�ыhf�B�P�M�QV�ҡhf�H�A�U�R�Ћhf�Q�Bx��W�M����E��t�E ��t�hf�Q�J�E�P����у���t�hf�B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�hf���   P�BH�Ћhf�Q���ȋBxW�Ѕ�t"�M�Q�U�R�M���/  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��S/  �EP�M�Q�M�u��u�/  ����   �u���E���tA��t<��uZ�hf���   �M�PHQ�ҋhf�Q���ȋBxV�Ѕ�u-�   ^��]Ëhf���   �E�JTP��VP�[�������uӍUR�E�P�M��/  ��u�3�^��]����������V��~ u>���t�hf�Q<P�B�Ѓ��    W�~��t���ʞ��W��������F    _^��������U��E�M�UP��P�EjP������]��������������̸   �����������U��V�u��t���u6�EjP��������u3�^]Ë�������t���t��U3�;P��I#�^]������̡hf�H\�������U��hf�H\�AV�u�R�Ѓ��    ^]�������������̡hf�P\�BQ�Ѓ���������������̡hf�P\�BQ�Ѓ����������������U��hf�P\�EPQ�J�у�]� ����U��hf�P\�EP�EPQ�J�у�]� U��hf�P\�EPQ�J�у�]� ���̡hf�P\�BQ�Ѓ����������������U��hf�P\�EPQ�J �у�]� ����U��hf�P\�EP�EPQ�J$�у�]� U��hf�P\�EP�EP�EPQ�J(�у�]� ������������U��hf�P\�EPQ�J0�у�]� ����U��hf�P\�EPQ�J@�у�]� ����U��hf�P\�EPQ�JD�у�]� ����U��hf�P\�EPQ�JH�у�]� ���̡hf�P\�B4Q�Ѓ����������������U��hf�P\�EP�EPQ�J8�у�]� U��hf�P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu��Ƶ���hf�H\�QV�҃���S��諵��3���~=��I �hf�H\�U�R�U��EP�A(VR�ЋM��Q���x����U�R���m���F;�|�_^[��]� ���������������U���VW�}�E��P��蘱���}� ��   �hf�Q\�BV�Ѓ��M�Q���q����E���t]S3ۅ�~H�I �UR���U����E�P���J����E;E�!���hf�Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U��V�u�F��F�����������������,0  ����������D�Ez��^��P�X]��������������N�X�N^�X]��������P�P�P�P �P(�P0�P8�P@�PH�PP�PX����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��5�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A��%����������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E������X�X]� ̋�3ɉ�H�H�H�V��V������FP����3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  S�]���q  ��؋�U��M�U�>�U��@�����@�U��@�B�@�������@���@�   ;����U��p  �w�����  �w�������F�B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]؋�R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ɍU��R�[�[������E��KH��P�E�SL��H�щKP�P�ST�H�KX�P�����S\��z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����M��}������3�3����u��u�|+�A�����B�4�u�0u��u�p�����u�u�U�E;�}�Q���E����U��U��1���@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���@�D��KX�@�U�����]��C���@�K0���@�KH���C ��C�@�K8���@�KP���C(��C�C@�H���@3����KX���U��r  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������]��E�E����]���E����]��E׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���@�   �KXE)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� ������������h�fPh_� � ������������������h�fjh_� ���������uË@����U��V�u�> t/h�fjh_� ���������t��U�M�@R�Ѓ��    ^]���U��Vh�fjh_� ����������t�@��t�MQ����^]� 3�^]� �������U��Vh�fjh_� ���Y�������t�@��t�MQ����^]� 3�^]� �������U��Vh�fjh_� ����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�fjh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh�fj h_� ����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh�fj$h_� ���I�������t�@$��t�MQ����^]� 2�^]� �������Vh�fj(h_� ����������t�@(��t��^��3�^������Vh�fj,h_� �����������t�@,��t��^��3�^������U��Vh�fj0h_� ����������t�@0��t�MQ����^]� 3�^]� �������U��Vh�fj4h_� ���i�������t�@4��t�M�UQR����^]� ���^]� ��Vh�fj8h_� ���,�������t�@8��t��^��3�^������U��Vh�fj<h_� �����������t�@<��t�MQ����^]� ��������������U��Vh�fj@h_� ����������t�@@��t�MQ����^]� ��������������U��Vh�fjDh_� ���y�������t�@D��t�MQ����^]� 3�^]� �������U��Vh�fjHh_� ���9�������t�@H��t�MQ����^]� ��������������Vh�fjLh_� �����������t�@L��t��^��3�^������Vh�fjPh_� �����������t�@P��t��^��3�^������Vh�fjTh_� ����������t�@T��t��^��^��������Vh�fjXh_� ���l�������t�@X��t��^��^��������Vh�fj\h_� ���<�������t�@\��t��^��^��������U��Vh�fj`h_� ���	�������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�fjdh_� �����������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh�fjhh_� ����������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh�fjlh_� ���9�������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�fjph_� �����������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh�fjth_� ����������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�fjxh_� ���i�������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh�fj|h_� ���)�������t�@|��t�MQ����^]� 3�^]� �������U��Vh�fh�   h_� �����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�fh�   h_� ����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�fh�   h_� ���6�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�fh�   h_� �����������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�fh�   h_� ����������t���   ��t�MQ����^]� 3�^]� �U��Vh�fh�   h_� ���F�������t���   ��t�MQ����^]� ��������U��Vh�fh�   h_� ����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�fh�   h_� ����������t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E����������m������U�_��^�U�[���U�������������������������  ����������D�Ez����P�X��]� �������E�����E����X�M��X��]� �����U���@�P&�A���E�    �����]��]��]��H&�������]��]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�q����F�@��R�M��_����~���Q�M��M����v;�t�v��P�M��7����M����m��M�u�_^[�M�UQR�M��������]� ��������������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$��-�E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��B-X-k--�-����U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�G����FP�>���3����F�F^��U��SV��WV�"����^S�����E3����~�~;�t_�hf�Q���   hX&��jIP�у��;�t9�}��t;�hf�B���   hX&��    jNQ�҃����uV������_^3�[]� �E�~_�F^�   []� ����������U��SV��WV�r����^S�i����}3Ƀ��N�N;���   9��   �G;���   �hf�Q���  hX&��jlP�у����t=� t@�G��t9�hf�JhX&��    ���  jqR�Ѓ����u������_^3�[]� �O�N�G�Q��    R�F�QP�  �����t�N�WP��QPR�x  ��_^�   []� ���������U��SV��WV�r����~W�i���3Ƀ��N�N9M��   �E;���   ��    �hf�H���  hX&h�   S�҃����t=�} tH�E��tA�hf�Q���  hX&��h�   P�у����u������_^3�[]� �U�V�,�F   �hf�H���  hX&h�   j�҃����t��E�M�F�PSPQ�q  �E����t!�V�?�W�RWP�U  ��_^�   []� ��M�_^�   []� ���U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��S�]V��3�W�~���F�F�CV;C��   贽��W讽��3��F�F�hf�Q���   hX&jIj�Ѓ������   �hf�Q���   hX&jNj�Ѓ����uV�V�����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� ����W�
���3��F�F�hf�B���   hX&jIj�у����t[�hf�B���   hX&jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP��������^]� ����������U��U��t�M��t�E��tPRQ�@  ��]������������U��E��u�E�M��f��f�   ]� �����������U��EHV����   �$��4�   ^]á�f@��f��uT�EP�����=�.  }�����^]Ëu��t�h�&jmh�fj�[�������t ���p����f��tV���t���   ^]���f    �   ^]ËM�UQR�U���������H^]�^]�p���-�fu.�"���m�����f��t���q��V��������f    �   ^]Ã��^]ÍI  4�4�4�3�4~4U��hf���   �BXQ�Ѓ���u]� �hf�Q|�M�RQ�MQP�҃�]� ���U��hf���   �BXQ�Ѓ���u]� �hf�Q|�M�R8Q�MQP�҃�]� ���U��EV��j ��hf�Qj j P�B�ЉF����^]� ��̡hfVj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� �hf�Q�MP�EP�Q�JP�у��F�   ^]� �N��Q��Q E��Q�D��Q�D��QVD��Q��Q�M��QrD��Q�C��QaCË�U�������;  �} ��ft��  ��]�; Qu���A  ��U��EVW��u|P�*  Y��u3��  �  ��u�*  ���*  � �Ԃ��(  ��f��"  ��}�  ����'  ��| �}%  ��|j �   Y��u��f�   �%  ��3�;�u19=�f~���f9=,ju�;"  9}u{��$  �  �*  �j��uY�q  h  j�  ��YY;��6���V�5�Q�5�i��  Y�Ѕ�tWV�  YY� �N���V�  Y�������uW�,  Y3�@_^]� jh�D�+  ����]3�@�E��u9�f��   �e� ;�t��u.��&��tWVS�ЉE�}� ��   WVS�r����E����   WVS�a����E��u$��u WPS�M���Wj S�B�����&��tWj S�Ѕ�t��u&WVS�"�����u!E�}� t��&��tWVS�ЉE��E������E���E��	PQ�*  YYËe��E�����3���*  Ë�U��}u�s,  �u�M�U�����Y]� ���̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�Ë�Q��&��,  YË�U��V��������EtV����Y��^]� ����U��WV�u�M�}�����;�v;���  ��   r�=�� tWV����;�^_u^_]�"1  ��   u������r*��$�T;��Ǻ   ��r����$�h:�$�d;��$��:�x:�:�:#ъ��F�G�F���G������r���$�T;�I #ъ��F���G������r���$�T;�#ъ���������r���$�T;�I K;8;0;(; ;;;;�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�T;��d;l;x;�;�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��<�����$��<�I �Ǻ   ��r��+��$��;�$��<�<(<P<�F#шG��������r�����$��<�I �F#шG�F���G������r�����$��<��F#шG�F�G�F���G�������V�������$��<�I �<�<�<�<�<�<�<�<�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��<�� ===,=�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̺PQ�!0  �PQ�/  �Ƀ=�ft�����=  �����z�����������������̃=�� �D  ���\$�D$%�  =�  u�<$f�$f��f���d$��C  � �~D$f('f(�f(�fs�4f~�fT@'f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�@  ���D$��~D$f��f(�f��=�  |!=2  �fT '�\�f�L$�D$����f�0'fV0'fT 'f�\$�D$�jh E�$  �e� �u;5��w"j�E  Y�e� V�$M  Y�E��E������	   �E��$  �j�D  YË�U��V�u�����   SW�= �=Dk u�R+  j�)  h�   �*  YY�����u��t���3�@P���uV�S���Y��u��uF�����Vj �5Dk�׋؅�u.j^9�ot�u��O  Y��t�u�{����O  �0�~O  �0_��[�V��O  Y�jO  �    3�^]������̋T$�L$��ti3��D$��u��   r�=�� t�P  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh E�#  �u��tu�=��uCj�C  Y�e� V�C  Y�E��t	VP��C  YY�E������   �}� u7�u�
j�oB  Y�Vj �5Dk� ��u�hN  ��� P�N  �Y��"  Ë�U��QSVW�5Ȃ�  �5Ă���}��t  ��YY;���   ��+ߍC��rwW�uO  ���CY;�sH�   ;�s���;�rP�u��S  YY��u�G;�r@P�u��=  YY��t1��P�4��  Y�Ȃ�u�  ���V�v  Y�Ă�EY�3�_^[�Ë�Vjj �  ��V�O  ���Ȃ�Ă��ujX^Ã& 3�^�jh@E�!  �  �e� �u�����Y�E��E������	   �E��!  ��  Ë�U���u���������YH]����������̃��$��O  �   ��ÍT$�O  R��<$�D$tQf�<$t�`O  �   �u���=�f ��O  �   ��Q��O  �  �u,��� u%�|$ u���5O  �"��� u�|$ u�%   �t����- S�   �=�f �vO  �   ��Q�N  ZË�U��EV���F ��uc��  �F�Hl��Hh�N�;8]t�T\�Hpu��Y  ��F;X[t�F�T\�Hpu�IR  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P��\  ��e�F�P�[  ��Yu��P�\  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P��[  �M��E��M��H��EP�\  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�s`  @PV�V��\  ��^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M�������3�;�u+��I  j_VVVVV�8�WY  ���}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�I  j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]hP'SV��_  ��3ۅ�tSSSSS�hW  ���N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�pt�90uj�APQ�u[  ���}� t�E��`p�3�_^[�Ë�U���,� Q3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�a  3ۃ�;�u�hH  SSSSS�0��W  �����o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q�$_  ��;�t���u�E�SP�u��V�u��������M�_^3�[�O����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �C���9}}�}�u;�u+�~G  j^WWWWW�0��V  ���}� t�E�`p����  9}vЋE��� 9Ew	�@G  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�J  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� ��_  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �y_  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�������u�E�8 u���} �4����$�p���WF�_  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP��]  0�F�U�����;�u��|��drj jdRP�]  0��U�F����;�u��|��
rj j
RP�]  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N�������u-�D  j^�03�PPPPP�S  ���}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V�������}� t�E��`p�3�_^[�Ë�U���,� Q3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�[  3ۃ�;�u�C  SSSSS�0�uR  �����Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P��Y  ��;�t���u�E�SV�u���`������M�_^3�[�
����Ë�U���0� Q3ŉE��ESV�uWj_W�M�Q�M�Q�p�0��Z  3ۃ�;�u�SB  SSSSS�8�Q  �����   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW�$Y  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[�����Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3����Q�6�  ��Y���(r�_^Ë�Vh   h   3�V��Z  ����tVVVVV��N  ��^Ë�U����`'�]��X'�]��E��u��M��m��]����]�����z3�@��3���h�'� ��thh'P� ��tj ���������U���(  ��g��g��g��g�5�g�=�gf��gf��gf��gf��gf�%�gf�-�g���g�E ��g�E��g�E��g������� g  ��g��f��f	 ���f   � Q�������$Q�������0 �gj�Z  Yj �, h�'�( �=g uj��Y  Yh	 ��$ P�  �Ë�U��V�5�Q�58 �օ�t!��Q���tP�5�Q���Ѕ�t���  �'��'V�4 ��uV�  Y��th�'P� ��t�u�ЉE�E^]�j ����YË�U��V�5�Q�58 �օ�t!��Q���tP�5�Q���Ѕ�t���  �'��'V�4 ��uV�   Y��th�'P� ��t�u�ЉE�E^]��< � ��V�5�Q�8 ����u�5�i�e���Y��V�5�Q�@ ��^á�Q���tP�5�i�;���Y�Ѓ�Q���Q���tP�D ��Q��c1  jh`E�  ��'V�4 ��uV�a  Y�E�u�F\((3�G�~��t$h�'P� �Ӊ��  h�'�u��Ӊ��  �~pƆ�   CƆK  C�Fh0Wj�2  Y�e� �vh�H �E������>   j��1  Y�}��E�Fl��u�8]�Fl�vl�qI  Y�E������   �  �3�G�uj��0  Y�j��0  YË�VW� �5�Q�������Ћ���uNh  j��  ��YY��t:V�5�Q�5�i�����Y�Ѕ�tj V�����YY� �N���	V����Y3�W�L _��^Ë�V��������uj�>  Y��^�jh�E�  �u����   �F$��tP�P���Y�F,��tP�B���Y�F4��tP�4���Y�F<��tP�&���Y�F@��tP����Y�FD��tP�
���Y�FH��tP�����Y�F\=((tP�����Yj�0  Y�e� �~h��tW�P ��u��0WtW����Y�E������W   j�P0  Y�E�   �~l��t#W�cH  Y;=8]t��`\t�? uW�oF  Y�E������   V�f���Y��  � �uj�/  YËuj�/  YË�U��=�Q�tK�} u'V�5�Q�58 �օ�t�5�Q�5�Q���ЉE^j �5�Q�5�i����Y���u�x�����Q���t	j P�@ ]Ë�VW��'V�4 ��uV�R  Y�����^  �5 h�'W��h�'W��i��h�'W��i��h�'W��i�փ=�i �5@ ��it�=�i t�=�i t��u$�8 ��i�D ��i�P�5�i��i�< ��Q�����   �5�iP�օ���   �_  �5�i�����5�i��i�����5�i��i�����5�i��i�u�������i��,  ��teh�R�5�i�����Y�У�Q���tHh  j�   ��YY��t4V�5�Q�5�i����Y�Ѕ�tj V�y���YY� �N��3�@��$���3�_^Ë�U��VW3��u�������Y��u'9�ivV�T ���  ;�iv��������uʋ�_^]Ë�U��VW3�j �u�u�qS  ������u'9�ivV�T ���  ;�iv��������uË�_^]Ë�U��VW3��u�u�ET  ��YY��u,9Et'9�ivV�T ���  ;�iv��������u���_^]Ë�U��W��  W�T �u�4 ���  ��`�  w��t�_]Ë�U���a  �u�  �5�Q�D���h�   �Ѓ�]Ë�U��h(�4 ��th (P� ��t�u��]Ë�U���u�����Y�u�X �j�n,  Y�j�+  YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=�& th�&�U  Y��t
�u��&Y�B���hD!h,!����YY��uBh$a������ !�$(!�c����=Ђ YthЂ�bU  Y��tj jj �Ђ3�]�jh�E�  j�+  Y�e� 3�C90j��   �,j�E�(j�} ��   �5Ȃ�����Y���}؅�tx�5Ă����Y���u܉}�u����u�;�rW����9t�;�rJ�6��������������5Ȃ�~������5Ă�q�����9}�u9E�t�}�}؉E����u܋}��hT!�H!�_���Yh\!�X!�O���Y�E������   �} u(�0jj�)  Y�u�����3�C�} tj�)  Y��7
  Ë�U��j j�u�������]�jj j ������Ë�V������V�5  V�W  V�C  V��  V��V  V��T  V�  V�T  hY������$��Q^�jTh�E�r	  3��}��E�P�h �E�����j@j ^V�&���YY;��  ����5����   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@�����   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M��������� ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=��|���=���e� ��~m�E����tV���tQ��tK�uQ�d ��t<�u���������4����E� ���Fh�  �FP�mU  YY����   �F�E�C�E�9}�|�3ۋ���5������t���t�N��r�F���uj�X�
��H������P�` �����tC��t?W�d ��t4�>%�   ��u�N@�	��u�Nh�  �FP��T  YY��t7�F�
�N@�����C���g����5���\ 3��3�@Ëe��E���������p  Ë�VW����>��t1��   �� t
�GP�l ���@   ;�r��6������& Y������|�_^Ã=̂ u�=  V�5�fW3���u����   <=tGV�H  Y�t���u�jGW�n�����YY�=j��tˋ5�fS�BV�\H  ��C�>=Yt1jS�@���YY���tNVSP��H  ����t3�PPPPP�L@  �����> u��5�f�
����%�f �' ���   3�Y[_^��5j������%j ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�S  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#��R  Y��t��M�E�F��M��E���R  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9̂u��:  h  �8jVS�<k�p �Ԃ�5 j;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�q�����Y;�t)�U��E�P�WV�}�������E���H�j�5j3�����_^[�Ë�U��@k��SV�5� W3�3�;�u.�֋�;�t�@k   �#� ��xu
jX�@k��@k����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5� SSS+�S��@PWSS�E��։E�;�t/P����Y�E�;�t!SS�u�P�u�WSS�օ�u�u�����Y�]��]�W�| ���\��t;�u��x ��;��r���8t
@8u�@8u�+�@P�E��0�����Y;�uV�t �E����u�VW�������V�t ��_^[�Ë�V��D��DW��;�s���t�Ѓ�;�r�_^Ë�V��D��DW��;�s���t�Ѓ�;�r�_^Ë�U��3�9Ej ��h   P�� �Dk��u]�3�@���]Ã=��uWS3�9��W�= ~3V�5����h �  j �v��� �6j �5Dk�׃�C;��|�^�5��j �5Dk��_[�5Dk�� �%Dk �Ë�U��QQV�G��������F  �V\�0RW�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   �$R�=(R���;�}$k��~\�d9 �=$R�(RB߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]��h�cd�5    �D$�l$�l$+�SVW� Q1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35 QW��E� �E�   �{���t�N�38�����N�F�38�����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���8N  �E���|@G�E��؃��u΀}� t$����t�N�38�����N�V�3:�����E�_^[��]��E�    �ɋM�9csm�u)�=�� t h����H  ����t�UjR������M��M  �E9Xth QW�Ӌ���M  �E�M��H����t�N�38�����N�V�3:�p����E��H���qM  �����9S�R���h QW���M  ������U���� Q�e� �e� SW�N�@��  ��;�t��t	�У$Q�`V�E�P�� �u�3u��� 3�� 3��� 3��E�P�� �E�3E�3�;�u�O�@����u������5 Q�։5$Q^_[��jh�E�r����e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E��t���Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[���������3��jhF����j�,  Y�e� �u�N��t/�Lk�Hk�E��t9u,�H�JP�V���Y�v�M���Y�f �E������
   ����Ë���j��  Y���������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�U���(  � Q3ŉE��@RVtj
��   Y�G  ��tj�G  Y�@R��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P�I�������������(�����0���j ǅ����  @��������,����, ��(���P�( j����̋�U��QQS�]VW3�3��}�;�HRt	G�}���r���w  j�L  Y���4  j�sL  Y��u�=�f�  ���   �A  hH.�  S�PkW�<  ����tVVVVV�4  ��h  �ikVj �ml �p ��u&h0.h�  V�O<  ����t3�PPPPP��3  ��V�;  @Y��<v8V�;  ��;�j�dnh,.+�QP�K  ����t3�VVVVV�3  ���3�h(.SW�kJ  ����tVVVVV�n3  ���E��4�LRSW�FJ  ����tVVVVV�I3  ��h  h .W�H  ���2j��` ��;�t$���tj �E�P�4�LR�6��:  YP�6S�� _^[��j�K  Y��tj��J  Y��u�=�fuh�   �)���h�   ����YYË�U��E�ln]�U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ë�U��� S3�9]u ��"  SSSSS�    �K2  ������   �MV�u;�t!;�u�"  SSSSS�    �2  ������S�����E�;�w�M�W�u�E��u�E�B   �u�u�P�u��GK  ����;�t�M�x�E����E�PS�I  YY��_^[�Ë�U���uj �u�u�u�5�����]�����U���0���S�ٽ\�����=X] t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=X] t�#  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����,  �   [�À�8�����=�f uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ��.�����������x.����s4��.�,ǅr���   ��.�����������p.����v��.VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�T  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����D   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Àzuf��\���������?�f�?f��^���٭^����S�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����S�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����S���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������- S��p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t�������0S u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t�@S���@S���l$����DS���DS���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r �������HS�|$�l$�ɛ�l$������l$��Ã�,��?�$��S����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  ������LS �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����|S�Ƀ�u�\$0�|$(���l$�-�S�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�lS�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���dS�|$�dS�<$� �|$$�D$$   �D$(�l$(���dS�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  ������LS �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����|S�Ƀ�u�\$0�|$(���l$�-�S�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�lS�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���dS�|$�dS�<$� �|$$�D$$   �D$(�l$(���dS�<$�l$$�Q�����0Z�����0Z�������@���������Ë�U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9pnt�5���T���Y�����M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E�\/��M��]�Q��]���]���Y����  �z  � "   �  �E�X/��M��]�Q��E�   �]���]���Y�j  �E�   �E�X/��E�P/��]���]���"  �M��E�P/�r����E�L/�׉M��E�L/�Z����E�\/놃�tNIt?It0It ��t����   �E�D/��E�</��E�\/����E�\/�x����E�   ��������   �E�   �E�4/��������������   �$�W��E�L/��E�P/��E�X/��E�,/��E�$/��E�/�y����E�/�m����E�/��E�/��E�/��M����]���]�M��]�Q�E�   ��Y��u��  � !   �E��_^[�þ�ǀЀـ��v���`�W�����%�� �������3�Ë�U��QQSV���  V�5�T�K  �EYY�M�ظ�  #�QQ�$f;�uU�?J  YY��~-��~��u#�ESQQ�$j��H  ���rVS�MK  �EYY�d�ES��!���\$�E�$jj�?�I  �]��EY�]�Y����DzVS�K  �E�YY�"�� u��E�S���\$�E�$jj�H  ��^[�Ë�VW3��xn�<��Tu���T�8h�  �0���6.  YY��tF��$|�3�@_^Ã$��T 3����S�l V��TW�>��t�~tW��W�f����& Y�����U|ܾ�T_���t	�~uP�Ӄ����U|�^[Ë�U��E�4ŘT�� ]�jh0F�7���3�G�}�3�9Dku�,���j�z���h�   ����YY�u�4��T9t���nj����Y��;�u�  �    3��Qj
�Y   Y�]�9u,h�  W�--  YY��uW蔼��Y�m  �    �]���>�W�y���Y�E������	   �E�������j
�(���YË�U��EV�4ŘT�> uP�"���Y��uj�����Y�6�� ^]Ë�U�������k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   ��o����   ����5� h @  ��H� �  SQ�֋����o�   ���	P��o�@�������    ��o�@�HC��o�H�yC u	�`���o�x�ueSj �p�֡�o�pj �5Dk� �����ok����+ȍL�Q�HQP�  �E�����;�ov�m�������E��o�=��[_^�á��V�5��W3�;�u4��k�P�5��W�5Dk�� ;�u3��x����5�����k�5��h�A  j�5Dk� �F;�t�jh    h   W�� �F;�u�vW�5Dk� 뛃N��>�~����F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�� ��u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U�������Mk���������M���SI�� VW}�����M���������3���U��������S�;#U�#��u
���];�r�;�u�����S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1����	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t����C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;�ou�M�;��u�%�o �M���B_^[�Ë�U��E3�;͸UtA��-r�H��wjX]ËͼU]�D���jY;��#���]�������u� WÃ��������u�$WÃ�Ë�U��V������MQ�����Y�������0^]Ë�U��E��o]Ë�U���5�o�����Y��t�u��Y��t3�@]�3�]�U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jhPF�����3��]3�;���;�u�y����    WWWWW��  ������S�=��u8j����Y�}�S�A���Y�E�;�t�s���	�u���u��E������%   9}�uSW�5Dk�� ���������3��]�u�j�����Y���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�2  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��`/�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z���/�����������|/�����   s���/���/�����������t/�����   v���/�����U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�-���3��ȋ��~�~�~����~����0W���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  � Q3ŉE�SW������P�v�� �   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R�j�����C�C��u�j �v�������vPW������Pjj �X?  3�S�v������WPW������PW�vS�9=  ��DS�v������WPW������Ph   �vS�=  ��$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[������jhpF������(������T\�Gpt�l t�wh��uj �[���Y��������j�,���Y�e� �wh�u�;5X[t6��tV�P ��u��0WtV�V���Y�X[�Gh�5X[�u�V�H �E������   뎋u�j�����YË�U���S3�S�M�蟬����o���u��o   �� 8]�tE�M��ap��<���u��o   �� �ۃ��u�E��@��o   ��8]�t�E��`p���[�Ë�U��� � Q3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�`[��   �E��0=�   r����  �p  ����  �d  ��P�� ���R  �E�PW�� ���3  h  �CVP芨��3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�C����M��k�0�u���p[�u��*�F��t(�>����E���\[D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C��d[Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95�o�X�������M�_^3�[������jh�F������M���������}�������_h�u�u����E;C�W  h   �8���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�P ��u�Fh=0WtP�2���Y�^hS�=H ���Fp��   �T\��   j����Y�e� �C��o�C��o�C��o3��E��}f�LCf�E�o@��3��E�=  }�L��PY@��3��E�=   }��  ��XZ@���5X[�P ��u�X[=0WtP�y���Y�X[S���E������   �0j�&���Y��%���u ��0WtS�C���Y�����    ��e� �E�����Ã=̂ uj��V���Y�̂   3�Ë�U��SV�u���   3�W;�to=X_th���   ;�t^9uZ���   ;�t9uP�ʥ�����   �z;  YY���   ;�t9uP詥�����   �;  YY���   葥�����   膥��YY���   ;�tD9u@���   -�   P�e������   ��   +�P�R������   +�P�D������   �9��������   �=�^t9��   uP��8  �7����YY�~P�E   ��X\t�;�t9uP����Y9_�t�G;�t9uP�֤��Y���Mu�V�Ǥ��Y_^[]Ë�U��SV�5H W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�X\t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5P W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�X\t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Å�t7��t3V�0;�t(W�8�����Y��tV�E����> Yu��`\tV�Y���Y��^�3��jh�F�u���輵����T\�Fpt"�~l t襵���pl��uj ����Y�������j����Y�e� �Fl�=8]�i����E��E������   ��j����Y�u�Ë�U��E�p]Ë�U���(  � Q3ŉE������� SjL������j P�/�����������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������0 j ���, ��(���P�( ��u��uj�H  Yh ��$ P�  �M�3�[�����Ë�U���5p�ı��Y��t]��j�	  Y]������U����u�M������E����   ~�E�Pj�u�A8  ������   �M�H���}� t�M��ap��Ë�U��=�o u�E�(]�A��]�j �u����YY]Ë�U���SV�u�M�脣���]�   ;�sT�M胹�   ~�E�PjS�7  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�8  YY��t�Ej�E��]��E� Y��1���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P��1  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=�o u�E�H���w�� ]�j �u�����YY]Ë�U���(� Q3ŉE�SV�uW�u�}�M��2����E�P3�SSSSW�E�P�E�P��A  �E�E�VP�f7  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�w����Ë�U���(� Q3ŉE�SV�uW�u�}�M�芡���E�P3�SSSSW�E�P�E�P�SA  �E�E�VP�<  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�ϔ������������������U��WV�u�M�}�����;�v;���  ��   r�=�� tWV����;�^_u^_]�"�����   u������r*��$�T���Ǻ   ��r����$�h��$�d���$���x���Ȣ#ъ��F�G�F���G������r���$�T��I #ъ��F���G������r���$�T��#ъ���������r���$�T��I K�8�0�(� �����D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�T���d�l�x����E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�������$����I �Ǻ   ��r��+��$����$����(�P��F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ��������Ĥ̤Ԥ��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$���� ���,��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��MS3�VW;�t�};�w�1���j^�0SSSSS���������0�u;�u��ڋъ�BF:�tOu�;�u������j"Y�����3�_^[]Ë�U��MSV�u3�W�y;�u�����j^�0SSSSS�.��������   9]v݋U;ӈ~���3�@9Ew����j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�a���@PWV�������3�_^[]Ë�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���H���u��P������Ɂ���  �P���t�M�_^f�H[�Ë�U���0� Q3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��A  �uЉC�E։�EԉC�E�P�uV������$��t3�PPPPP�<������M�_�s^��3�[�R������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j蹭��YË�U��E�M%����#�V������t1W�}3�;�tVV�J  YY�����j_VVVVV�8� �������_��uP�u��t	�QJ  ���HJ  YY3�^]Ã%�� �jh�F蘹���M3�;�v.j�X3���;E�@u�4����    WWWWW������3���   �M��u;�u3�F3ۉ]���wi�=��uK������u�E;��w7j����Y�}��u����Y�E��E������_   �]�;�t�uWS�V�����;�uaVj�5Dk� ��;�uL9=�ot3V�����Y���r����E;��P����    �E���3��uj�G���Y�;�u�E;�t�    ���̸���jh�F�z����]��u�u�����Y��  �u��uS�2���Y�  �=����  3��}�����  j����Y�}�S�����Y�E�;���   ;5��wIVSP��������t�]��5V����Y�E�;�t'�C�H;�r��PS�u��L���S�����E�SP������9}�uH;�u3�F�u������uVW�5Dk� �E�;�t �C�H;�r��PS�u������S�u��b������E������.   �}� u1��uF������uVSj �5Dk�� ����u�]j�����YË}����   9=�ot,V�1���Y������������9}�ul��� P�v���Y��_����   ����9}�th�    �q��uFVSj �5Dk�� ����uV9�ot4V�����Y��t���v�V����Y�Z����    3��ٶ����G����|�����u�9������ P������Y��������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�hGh�cd�    P��SVW� Q1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh0G�����N����@x��t�e� ���3�@Ëe��E������(���� ����h]��U���Y�pË�U��E� p�$p�(p�,p]Ë�U��E�0RV9Pt��k�u��;�r�k�M^;�s9Pt3�]��5(p�i���Y�j hPG�[���3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�������}؅�u����a  � p� p�`�w\���]���������Z�Ã�t<��t+Ht�����    3�PPPPP������뮾(p�(p��$p�$p�
�,p�,p�E�   P襠���E�Y3��}���   9E�uj蘩��9E�tP�����Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.�$R�M܋(R�$R�9M�}�M�k��W\�D�E���������E������   ��u�wdS�U�Y��]�}؃}� tj ����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3������Ë�U��E�4p]Ë�U��E�8p]�jhpG荲���e� �u�u�� �E��/�E� � �E�3�=  �����Ëe�}�  �uj�L �e� �E������E�����Ë�U����u�M�萑���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]���SVW�T$�D$�L$URPQQh4�d�5    � Q3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�F  �   �C�$F  �d�    ��_^[ËL$�A   �   t3�D$�H3��K���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�oE  3�3�3�3�3���U��SVWj j h۲Q�e  _^[]�U�l$RQ�t$������]� ��U���SVW�`����e� �=xp ����   h�7�� �����*  �5 h�7W�օ��  P誜���$�7W�xp��P蕜���$|7W�|p��P耜���$`7W��p��P�k���Y��p��thH7W��P�S���Y��p��p;�tO9�ptGP豜���5�p��褜��YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9�|p;�t0P�a���Y��t%�ЉE���t��p;�tP�D���Y��t�u��ЉE��5xp�,���Y��t�u�u�u�u����3�_^[�Ë�U��ES3�VW;�t�};�w����j^�0SSSSS���������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��e���j"Y����3�_^[]Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w�#���j^�0SSSSS����������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x��������j"Y���낋�U��MV3�;�|��~��u��f�(��f��f��n���VVVVV�    ����������^]Ë�U��E��t���8��  uP�Y���Y]Ë�U��QV�uV�wO  �E�FY��u����� 	   �N ����/  �@t������ "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�TM  �� ;�t�HM  ��@;�u�u��L  Y��uV�L  Y�F  W��   �F�>�H��N+�I;��N~WP�u�uK  ���E��M�� �F����y�M���t���t����������������Q�@ tjSSQ��B  #����t%�F�M��3�GW�EP�u�K  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u�C����8*u�ϰ?�d����} �^[]Ë�U���x  � Q3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������u�����u5�����    3�PPPPP������������ t
�������`p������
  �F@u^V��L  Y��Q���t���t�ȃ��������������A$u����t���t�ȃ������������@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw�����7��3��3�3�����7j��Y������;���	  �$�v���������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�������Q  Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u�T]������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P��I  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  �P]������P����Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7���������{G  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V�+���������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5�Q�$���Y�Ћ���������   t 9�����u������PS�5�Q�����Y��YY������gu;�u������PS�5�Q�А��Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�I7  ��0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u�P]�������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF�D  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t�������*}�������� Y���������������t������������������������� t
�������`p��������M�_^3�[�,s���Ð�������\�g���ۻ��S��QQ�����U�k�l$���   � Q3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�(  ��h��  ��x����  �>YYt�=X] uV�    Y��u�6��  Y�M�_3�^��q����]��[�3�Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u�� �M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M����X^��{L�H��M�����{,�X^�2��M�����z�X^���M�����z�H^��H^��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E����!�S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�X���� "   ]��K���� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���`];Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�U�������uV�,���Y�E�^�Ë�d]�h��  �u(�  �u�����E ���Ë�U��=X] u(�u�E���\$���\$�E�$�uj�/�����$]��4���h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   � Q3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=X] u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3���j����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-p^�]���t����-p^�]�������t
�-|^�]����t	�������؛�� t���]����jh�G葕��3�9��tV�E@tH9�^t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�^ �e��U�E�������e��U�q���Ë�U���� Q3ŉE�SV3�W��9�pu8SS3�GWh�8h   S�� ��t�=�p�� ��xu
��p   9]~"�M�EI8t@;�u�����E+�H;E}@�E��p����  ;���  ����  �]�9] u��@�E �5� 3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�*  ��;�t� ��  �P�o��Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5� SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�B)  ��;�tj���  ���P��n��Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�� ��t"SS9]uSS��u�u�u�VS�u �� �E�V�g���Y�u��^����E�Y�Y  �]�]�9]u��@�E9] u��@�E �u�6  Y�E���u3��!  ;E ��   SS�MQ�uP�u ��6  ���E�;�tԋ5� SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�,(  ��;�t����  ���P��m��Y;�t	� ��  �����3�;�t��u�SW�n�����u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��6  ���u������#u�W�<���Y��u�u�u�u�u�u�� ��9]�t	�u��n��Y�E�;�t9EtP�un��Y�ƍe�_^[�M�3��d���Ë�U����u�M���p���u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap��Ë�U��QQ� Q3ŉE���pSV3�W��;�u:�E�P3�FVh�8V�� ��t�5�p�4� ��xu
jX��p���p����   ;���   ����   �]�9]u��@�E�5� 3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�E&  ��;�t� ��  �P��k��Y;�t	� ��  ���؅�ti�?Pj S�l����WS�u�uj�u�օ�t�uPS�u�� �E�S�x����E�Y�u3�9]u��@�E9]u��@�E�u��3  Y���u3��G;EtSS�MQ�uP�u��3  ����;�t܉u�u�u�u�u�u�� ��;�tV�vl��Y�Ǎe�_^[�M�3��b���Ë�U����u�M���n���u$�M��u �u�u�u�u�u�������}� t�M��ap��Ë�U��V�u����  �v�l���v��k���v��k���v��k���v��k���v��k���6��k���v ��k���v$��k���v(�k���v,�k���v0�k���v4�k���v�k���v8�k���v<�k����@�v@�k���vD�|k���vH�tk���vL�lk���vP�dk���vT�\k���vX�Tk���v\�Lk���v`�Dk���vd�<k���vh�4k���vl�,k���vp�$k���vt�k���vx�k���v|�k����@���   ��j�����   ��j�����   ��j�����   ��j�����   ��j�����   ��j�����   �j�����   �j�����   �j�����   �j�����   �j����,^]Ë�U��V�u��t5�;X_tP�mj��Y�F;\_tP�[j��Y�v;5`_tV�Ij��Y^]Ë�U��V�u��t~�F;d_tP�'j��Y�F;h_tP�j��Y�F;l_tP�j��Y�F;p_tP��i��Y�F;t_tP��i��Y�F ;x_tP��i��Y�v$;5|_tV�i��Y^]��������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U���S�u�M��k���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�/����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M���j���E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�_N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC��_��+�_;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�_N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���_A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�_��_��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硠_��_�3�@�   ��_�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�_��M���Ɂ�   �ً�_]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�_N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC��_��+�_;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�_N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���_A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�_��_��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硸_��_�3�@�   ��_�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�_��M���Ɂ�   �ً�_]���@u�M�U�Y��
�� u�M�_[�Ë�U���|� Q3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u����SSSSS�    聻����3��N  �U�U��< t<	t<
t<uB��0�B���/  �$����Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�a#  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �"  =�����.  �c��`�E�;���  }�عpd�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��K
3��E��EԉE؉E܋E΋��  3�#�#ʁ� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uB�E����u9u�u9u�u3�f�E���  f;�u!B�C���u9su93u�ủuȉu���  �u��}��E�   �E��M���M���~R�DĉE��C�E��E��M��	� �e� ���O��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?�����  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋M��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9M�w�Mԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�B�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�U�f�EċE؉EƋE܉E�f�U��3�f�����e� H%   � ���e� �Ẽ}� �<����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[�M���ÐU�����2�w������	���}�,���U���t� Q3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�f��t�C-��C �u�}�f��u/��u+��u'3�f;�����$ f��C�C�C0�S3�@�  ��  f;���   3�@f��   �;�u��t��   @uh�A�Qf��t��   �u��u;h�A�;�u0��u,h�A�CjP������3���tVVVVV蔲�����C�*h�A�CjP������3���tVVVVV�h������C3��q  �ʋ�i�M  �������Ck�M��������3���f�M�c�ۃ�`�E�f�U�u�}�M�����  }�pd�ۃ�`�E�����  �E�T�˃������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE��P
3ɉM��M��M�M��M��3�� �  �u���  #�#֍4
����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��{����M�����?  ��  f;���  �E�3҉U��U��U�U��U��ɋ�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��V���3�3�f9u���H%   � ���E��\���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �^�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[�D���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95����  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��{���Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��U��SVWUj j h,��u�b!  ]_^[��]ËL$�A   �   t2�D$�H�3��K?��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h4�d�5    � Q3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y4�u�Q�R9Qu�   �SQ��_�SQ��_�L$�K�C�kUQPXY]Y[� ��������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ��U��j
j �u�  ��]�������Q�L$+ȃ����Y�*  Q�L$+ȃ����Y�  ��U��QQ�EV�u�E��EWV�E��  ���Y;�u蒕��� 	   �ǋ��J�u�M�Q�u�P�� �E�;�u� ��t	P脕��Y�ϋ������������D0� ��E��U�_^��jh�G�si������u܉u��E���u�)����  ����� 	   �Ƌ���   3�;�|;��r!������8����� 	   WWWWW�H������ȋ���������������L1��u&辔���8褔��� 	   WWWWW������������[P�  Y�}���D0t�u�u�u�u�������E܉U���V���� 	   �^����8�M���M���E������   �E܋U��h����u�@  YË�U���  �g  � Q3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�����0�ғ��VVVVV�    �5���������  SW�}�����4��������ǊX$�����(�����'�����t��u0�M����u&胓��3��0�g���VVVVV�    �ʢ�����C  �@ tjj j �u�~������u�i  Y����  ��D���  �V���@l3�9H�������P��4�� ����� ���`  3�9� ���t���P  �� ��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P�Z���Y��t:��4���+�M3�@;���  j��@���SP�[  �������  C��D����jS��@���P�7  �������  3�PPj�M�Qj��@���QP�����C��D����� �����\  j ��<���PV�E�P��(���� �4�� ���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4�� ����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@����D  Yf;�@����h  ��8����� ��� t)jXP��@����  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4�� ���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4�� ���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �� ��;���   j ��,���P��+�P��5����P��(���� �4�� ��t�,���;���� ��@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0�� ��t��,�����@��� ��8����� ��@�����8��� ul��@��� t-j^9�@���u�Z���� 	   �b����0�?��@����f���Y�1��(�����D@t��4����8u3��$�����    �"����  ������8���+�0���_[�M�3�^�d4����jh�G�'a���E���u�����  �ˌ��� 	   ����   3�;�|;��r!轌���8裌��� 	   WWWWW�������ɋ���������������L1��t�P��  Y�}���D0t�u�u�u�.������E���@���� 	   �H����8�M���E������	   �E��`����u�1  YË�U����ph   ��R��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u赋��� 	   3�]�V3�;�|;��r藋��VVVVV� 	   �������3���ȃ����������D��@^]ø�_á��Vj^��u�   �;�}�ƣ��jP�RR��YY�`q��ujV�5���9R��YY�`q��ujX^�3ҹ�_��`q��� ����`b|�j�^3ҹ�_W������������������t;�t��u�1�� B��P`|�_3�^��  �=(j t��  �5`q�;��YË�U��V�u��_;�r"��@bw��+�����Q�)���N �  Y�
�� V�� ^]Ë�U��E��}��P��~���E�H �  Y]ËE�� P�� ]Ë�U��E��_;�r=@bw�`���+�����P��}��Y]Ã� P�� ]Ë�U��M���E}�`�����Q�}��Y]Ã� P�� ]Ë�U��EV3�;�u蚉��VVVVV�    ������������@^]á Q��3�9�p����Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�$���j^SSSSS�0舘�������V�u�M��<���E�9X��   f�E��   f;�v6;�t;�vWSV�9�����ш��� *   �ƈ��� 8]�t�M��ap�_^[��;�t2;�w,覈��j"^SSSSS�0�
�����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�� ;�t9]�^����M;�t���� ��z�D���;��g���;��_���WSV�8�����O�����U��j �u�u�u�u�|�����]Ë�U���� Q3ŉE�j�E�Ph  �u�E� �� ��u����
�E�P����Y�M�3��/���Ë�U���4� Q3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5� �M�QP�֋� ��t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��4�����YF;�~[�����wS�D6=   w/������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�6��Y;�t	� ��  ���E���}�9}�t؍6PW�u��<7����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�� ��t`�]��[�� 9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�NM��YY�E�;�t+WWVPV�u�W�u��;�u�u��07��Y�}���}��t�MЉ�u�衬��Y�E��e�_^[�M�3��X-���Ë�U���� Q3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[�+���Ë�U���VW�u�M��7���E�u3�;�t�0;�u,����WWWWW�    �I������}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�����M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&�E����E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9�ouh@]�P������]����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ���U��MS3�;�VW|[;��sS������<����������@t5�8�t0�=�fu+�tItIuSj��Sj��Sj�� !���3������� 	   ��������_^[]Ë�U��E���u������  �ހ��� 	   ���]�V3�;�|";��s�ȃ�����������@u$踀���0螀��VVVVV� 	   ����������� ^]�jh�G�T���}����������4����E�   3�9^u6j
�u��Y�]�9^uh�  �FP����YY��u�]��F�E������0   9]�t�������������D8P�� �E��|T���3ۋ}j
��s��YË�U��E�ȃ����������DP�� ]Ë�U���� Q3ŉE�V3�95�etO�=Df�u�g  �Df���u���  �pV�M�Qj�MQP�!��ug�=�eu�� ��xuω5�eVVj�E�Pj�EPV�!P�� �Df���t�V�U�RP�E�PQ�!��t�f�E�M�3�^�y&������e   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��m2���E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�G���YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�� ���E�u�M;��   r 8^t���   8]��e����M��ap��Y����~��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�� ���:���뺋�U��j �u�u�u�������]�jhH��Q��3ۉ]�j�sr��Y�]�j_�}�;=��}W�����`q�9tD� �@�tP�  Y���t�E��|(�`q��� P�l �`q�4�p.��Y�`q�G��E������	   �E��Q���j�q��YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�C���YP�������;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�����P�  Y��Y��3�^]�jh0H�P��3��}�}�j�!q��Y�}�3��u�;5����   �`q��98t^� �@�tVPV�����YY3�B�U��`q���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u�`q�4�V�����YY��E������   �}�E�t�E��1P���j�o��Y�j����Y����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h<B�!�DfáDfV�5!���t���tP�֡@f���t���tP��^Ë�U��SV�uW3����;�u��z��WWWWW�    �&�������B�F�t7V�{���V����  V�����P�   ����}�����F;�t
P�+��Y�~�~��_^[]�jhXH�N���M��3��u3�;���;�u�@z���    WWWWW裉���������F@t�~�E��N���V����Y�}�V�*���Y�E��E������   �ՋuV�����Y�jhxH�$N���E���u��y��� 	   ����   3�;�|;��r�y��� 	   SSSSS�������Ћ����<�����������L��t�P�����Y�]���Dt1�u�g���YP�!��u� �E���]�9]�t�Ny���M��1y��� 	   �M���E������	   �E��M����u�)���YË�U��V�uWV� ���Y���tP�����u	���   u��u�@Dtj�����j�������YY;�tV�����YP�!��u
� ���3�V����������������Y�D0 ��tW�x��Y����3�_^]�jh�H�L���E���u�fx���  �Kx��� 	   ����   3�;�|;��r!�=x���8�#x��� 	   WWWWW膇�����ɋ���������������L1��t�P�g���Y�}���D0t�u�����Y�E����w��� 	   �M���E������	   �E��6L����u�����YË�U��V�u�F��t�t�v�(���f����3�Y��F�F^]�����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%� ������������h��U)��Y����̃=�f uK��f��t�hf�Q<P�B�Ѓ���f    ��f��tV�������V���������f    ^�                                                                                                                                                                                                                                                           �I J 0J BJ NJ ^J jJ |J �J �J �J �J �J K K (K 4K BK LK dK tK �K �K �K �K �K �K �K �K L ,L DL ^L tL �L �L �L �L �L �L �L M M 6M NM ^M lM xM �M �M �M �M �M �M �M N N $N :N JN \N nN �N �N �N �N �N �N �N �N O         �        �A�f��"��         }                9	0N       p   �B �0 bad allocation                    �?    USERNAME         @�@ikto    ikfrom  texturesearchpath   dst src fbx c4d c:\buildagent\work\b2b44f52c74c2f2a\src\source\convert.cpp  EXPORT_ERROR: An unknown error has occured  EXPORT_ERROR: An error occured while saving the document    EXPORT_ERROR: Destination bad format    EXPORT_ERROR: Source bad format EXPORT_ERROR: Source either does not exist or cannot be located EXPORT_ERROR: An error occured while loading the document   EXPORT_ERROR: FBX exporter not found    SUCCESS framerate=  version=    -UnityC4DFBXtmp -UnityC4DFBXout 0   Filtered:       Name: ' '   Plugin:     Processing  Scanning    -UnityC4DFBXcmd * (c) 2006-2011 Unity Technologies ApS - http://unity3d.com * Unity-C4DToFBXConverter for Cinema 4D R13. Version: 3.09  ����MbP?�C`� �m �C@�     c:\buildagent\work\b2b44f52c74c2f2a\sdk\r13\_api\c4d_baseobject.cpp c:\buildagent\work\b2b44f52c74c2f2a\sdk\r13\_api\c4d_general.h  %s     c:\buildagent\work\b2b44f52c74c2f2a\sdk\r13\_api\c4d_file.cpp       c:\buildagent\work\b2b44f52c74c2f2a\sdk\r13\_api\c4d_basetime.cpp             �? �Ngm��C   ����A  4&�k�  4&�kC(Dp� c:\buildagent\work\b2b44f52c74c2f2a\sdk\r13\_api\c4d_resource.cpp   #   M_EDITOR        �������������c:\buildagent\work\b2b44f52c74c2f2a\sdk\r13\_api\c4d_libs\lib_ngon.cpp  c:\buildagent\work\b2b44f52c74c2f2a\sdk\r13\_api\c4d_pmain.cpp  |6�a�a    pD�9              �?      �?3      3            �      0C       �       ��              e+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    �f gEncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:                �������             ��      �@      �              �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow       �?5�h!���>@�������             ��      �@      �            	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        �5�5�5�5�5�5t5l5`5T5�!�0|0h0H0,0L5D5(0@5<5854505,5 55555555 5�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4x4`4T4@4 4 4�3�3�3|3`3<33�2�2�2�2�2�2�2�2t2d2H2(2 2�1�1�1h1D1 1�0�0�0�!GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun 1#QNAN  1#INF   1#IND   1#SNAN  SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                            Q�D   RSDS3�����B��RTeFC�   C:\BuildAgent\work\b2b44f52c74c2f2a\src\obj\Unity-C4DToFBXConverter13_Win32_Release.pdb            pCxC    lP        ����    @   `C            �P�C           �C�C    �P        ����    @   �C            �P�C            DDxC    �P       ����    @   �C            �P<D           LDTD    �P        ����    @   <D            4Q�D           �D�D    4Q        ����    @   �D        �c 4� 4�                     ����    ����    �����8�8    ����    ����    ����    �>    ����    ����    ����    �@    ����    ����    ����    �A    ����    ����    ����    +R����    :R����    ����    ����    �S����    �S����    ����    ����    gY    ����    ����    ����/\3\    ����    ����    ����f+f    ����    ����    ����    g    ����    ����    ����    �    ����    ����    ����    !�    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    Y�    ����    ����    ����    ê    ����    ����    ����    (�    ����    ����    ����+�?�    ����    ����    ����}���    ����    ����    ����    w�    ����    ����    �������    ����    ����    ���� ��    ����    ����    ����     �    ����    ����    ����        ����    ����    ����    :    ����    ����    ����    �    ����    ����    ����    �        Q����    ����    ����    5    ����    ����    ����        ����    ����    ����    ��H         J                        �I J 0J BJ NJ ^J jJ |J �J �J �J �J �J K K (K 4K BK LK dK tK �K �K �K �K �K �K �K �K L ,L DL ^L tL �L �L �L �L �L �L �L M M 6M NM ^M lM xM �M �M �M �M �M �M �M N N $N :N JN \N nN �N �N �N �N �N �N �N �N O     ZGetTempPathA  KERNEL32.dll  �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �GetLastError  �HeapFree   GetProcAddress  �GetModuleHandleA  -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent �GetModuleHandleW  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �InterlockedIncrement  �SetLastError  �InterlockedDecrement  !Sleep ExitProcess �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA � DeleteCriticalSection �GetModuleFileNameA  JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW zWideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy WVirtualFree TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �WriteFile �LeaveCriticalSection  � EnterCriticalSection  TVirtualAlloc  �HeapReAlloc �HeapSize  [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �LoadLibraryA  �InitializeCriticalSectionAndSpinCount �RtlUnwind �GetLocaleInfoA  ZRaiseException  �LCMapStringA  MultiByteToWideChar �LCMapStringW  =GetStringTypeA  @GetStringTypeW  �SetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW x CreateFileA C CloseHandle AFlushFileBuffers              9	0N    RO          HO LO PO �3 pO   Unity-C4DToFBXConverter13.cdl c4d_main                                                                                                                                        |!    |!    B�     b�     a�     `�     ��    ��    qr            |!|!|!|!|!|!|!�&    .?AVGeSortAndSearch@@   �&    .?AVNeighbor@@  �&    .?AVDisjointNgonMesh@@  |!|!|!|!|!|!�&    .?AVBaseData@@  |!|!|!|!|!|!|!|!|!u�  s�  N�@���D        |!�&    .?AVtype_info@@     fmod         d=&q�p&q�p&q�p&q�p�p�p�p&q&q�p&qsqrt    O�O�O�O�O�O�O�O�O�O���������Y    �����
                                                                   x   
   |!                  �-   �-	   x-
   �,   �,   �,   `,   4,   �+   �+   �+   d+   <+   +   �*    �*!   �)"   �(x   �(y   �(z   �(�   �(�   �(       ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ���trzrr�r�r�r�r�r�r�r�r�r�r�r
ss.sNsSsmsrs�s�s�s�s�s�stt6tJtbtvt�t�t�t�t�t�tuu:u?uYu^u~u�u�u�u�u�u�uv"v6vNvbv�v�v�v�v�v�v�v  ?                                                                                                                                                                                                                                                                                                                         	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                                                                             abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     0W�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    �;����C                                                                                              X\            X\            X\            X\            X\                              X_        �90>�?�^`\   `\0W        �7�7�&         X/   \/   L/   P/   �8   �8!   �8   D/   </   ,/   �8   |8   /   /    /   $/   /   t8   /   l8   d8   \8   T8   L8"   H8#   D8$   @8%   88&   ,8      �      ���������              �       �D        � 0     �9�;    �A�A�A�A�A�A�A�A�A�A�A�A�A|AxAtApAlAhAdA`A\AXATAPALADA8A0A(AhA AAAA�@�@�@�@�@�@�@�@	         �^.   T_�p�p�p�p�p�p�p�p�pX_   .                 ���5      @   �  �   ����              �            �q    �q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �p     ����    PST                                                             PDT                                                             pb�b����        ����                 �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
       ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                             0"000A0N0d0�0�0�0�01'151D1t1�1�1�1�1�122�2�2�2b3�3�3�3444K4]4o4�4�4�4�4�4�4�45:5\5�5�56:6v6�6�6�67-7K7i7�7�7;8W8p8�8�89�9�9�9�9�9
:,:>:P:�:�:�:�:�:�:;!;3;?;N;g;�;�;�;�;�;�;
<<-<M<[<q<�<�<�<�<�<==*=J=d=x=�=�=�=�=�=>>e>�>�>�>�>�>9?�?�?�?      0  	040P0j0�0�0�0�0�011Q1�12w2�2�233\3n33�3�3�3�344/4X4j4|4�4�4�5�5�5�5�5�566-6A6V6k66�6�6�6�6�6�6%7,7L7j7�7�7�7�78#8=8T8e8w8�8�8�8�8�8�8�8�89$9b9�9�9:$:(:,:0:4:q:�:�:�:�:�:�:�:�:�:;";+;=;O;W;m;;�;�;�;<4<L<`<|<�<�<�<�<�<@=U=j=r=�=�=�=�=�=	>&>>>f>k>�>�>�>�>�>�>?#?8?J?\?e?{?�?�?�?�? 0  @  0 020;0Q0f0z0�0�0�0�0�0�0�01N1a1�1�1�1�1�1�1�124282<2@2D2H2L2P2T2X2\2`2�2�2�2�2�2�2�233(3M3a3w3�3�3�3�3�344$464V4r4�4�4�4�4�4�45!535E5V5h5z5�5�5�5�5 66$666G6Y6b6t6�6�6�6�6�677,7@7c7u7�7�7�7�7�7�78*8<8�8�8�8�8�809A9S9e9w9�9�9�9�9�9::T:t:�:�:�:�:�:;>;P;b;s;�;�;�;�;<7<A<=B=r=�=�=">U>�>�>%?5?u?�?   @  �   0:0�0�0�0E1�1�1�1%2u2�2353�3�3�3%4e4�4�45U5�5�5%6e6�6�6�67757�7�78B8�8�89b9�9�9:):3:`:e:�:�:�:;);e;�;�;�;E<i<�<�<�<&=O=�=�=�=>Y>�>�>�?�?�?�?�? P  �   040T0t0�0�0�0�0�0�01$1D1d1�1�1�1�12!2D2a2�2�2�2�2343T3t3�3�3�34!444T4t4�4�4�4�45/5T55�5�5�56-6<6a6t6�6�6�6�6�67T7t7�7�7�7848�8�8$9d9�9�9�9�9:$:D:d:�:�:�:�:$;D;t;�;�;�;<4<a<�<�<�<=1=T=�=�=�=>!>A>a>�>�>�>�>?!?A?a?�?�?�?�?   `  �   0$0T0t0�0�0�0141Q1t1�1�1�12D2t2�2�23R3q3�3�3�3�3$4Q4q4�4�4�4�4$5T5�5�5�5�5646d6�6�6�6�6�6!707T7�78A8T8t8�8�8�8!9A9q9�9�9�9:!:D:�:�:�:;4;d;�;�;�;:<{<�<�<�<=4=d=�=�=�=�=�=>J>d>�>�>?*?t?�?�?   p  �   r0�0!151J1m1�1�1�1#2F2o2�2�2�23X3�34T4d4�4�4�45C5W5u5�5�5�56$6T6t6�6�6�67$7q7�7�7�7818T8t8�8�8�849�9�9�9�9:O:n:�:�:�:;8;S;�;�;�;�;�;<6<f<�<�<�<�<�</=C=X=�=�=�=�=!>;>[>p>�>G?Z?�?�?�?�? �  �   0\0k2535�5�5�5�56T6o6$8(8,808k8p8�8�8�899D9t9�9�9�9:4:T:�:�:�:;4;T;t;�;�;�;�;<4<F<a<t<�<�<�<�<�<=4=q=�=�=�=�=>4>T>q>�>�>�>�>�>?$?D?d?�?�?�?�? �  �   040Q0d0�0�0�0�01$1t1�1�1�12$2D2d2�2�2�2�23$3d3�3�34c4�4�4545d5�5�5�5�5616A6T6t6�6�6�6�6)7=7�7�7�7�7$8D8d8�8�8�8�8929F9V9�9�9�9�9:$:P:d:t:�:�:�:;*;];k;~;�;�;�;�;�;<.<B<R<t<�<�<�<==E=s=�=�=�=�=�=>C>Y>g>v>�>�>�>?D?m?�?�?�?   �    0$0O0t0�0�0�0�0111D1d1�1�1�1�1242T2t2�2�2�2�2343Q3a3t3�3�3�3�34!4D4Y4k4�4�4�4�4�45$555C5d5u5�5�5�5�5�5�5646T6q6�6�6�6�6�67$7<7P7_7o7�7�7�7�7�7�7 8=8O8q8�8�8�8�8�89D9V9d9w9�9�9�9:4:Q:d:�:�:�:�:;$;D;d;�;�;�;�;�;�;<4<T<t<�<�<�<�<=4=T=n=�=�=�=�=�>??/?P?X?l?�?   �  (  0;0Q0u0�0�0�0141T1t1�1�1�1�1242Q2a2t2�2�2�2�2�2�2343S3a3p3�3�3�344!414A4Q4d4�4�4�4�4�4�45$5D5d5�5�5�5�56$6W6p6�6�6�6�6�67'797d7�7�7�7�78$8;8O8^8n8�8�8�8�8�8�89$9H9n9�9�9�9�9�9�9::4:R:f:u:�:�:�:;$;D;a;t;�;�;�;�;�;<4<T<t<�<�<�<�<=4=T=t=�=�=�=�=>4>T>t>�>�>�>�>$?P?t?�?�?�?�? �  �   040T0t0�0�0�0�0141T1t1�1�1�1�1242T2t2�2�2�2�23$3D3a3t3�3�3�3�3�34&4:4J4t4�4�4�4555R5D6d6~6�6�6�6�6?7a7�7�7�7�78$8T8f8�8�8�8�8$9D9a9�9�9�9�9:$:T:o:�:�:�:�:;$;T;�;�;�;�;<4<d<�<�<�<=$=Q=t=�=�=�=>4>T>t>�>�>�>�>?4?Q?d?�?�?�?�?   �  �   N0n0�0�0'1�1�12x2�2�283Z3}3�34&4�4�4�4S5|5�5�5�5D6�6747�7�78�8�8�8N9n9�9�9l:�:�:;q;�;�;<q<�<S=|=�=>>>S>�>�>?Q?g?�?   �  �   ,0�0�0�011$1T1t1�1�1�12$2a2�2�2�2�23$3W3�3�3�3�3.4G4[4z4�4�45!5D5a5�5�5>6C6H6M6o6�6�6�67747T7t7�7�7�7$8D8d8�8�8�8�8�89B9p9�9�9:@:n:�:�:�:;�;�;%<<<Q<Z<m<�<�<==Z=j=�=�=>>$>a>t>�>�>�>�>?!?4?T?|?�?�?�? �    $0D0a0�0�0I1e1�1�1I2e2�2�23,3H3d3�3�34%4�4�4!5�5�5�5�56$6J6X6g6�6�6�6'7[7�7�7�7�7�7
8$818>8V8i8{8�8�8�8�8�8�89(9D9U9h9�9�9�9�9�9�9�9::6:T:f:�:�:�:�:�:�:�: ;6;R;c;v;�;�;�;�;�;�;<<(<F<d<v<�<�<�<�<�<�<=0=F=b=t=�=�=�=�=�=>4>B>O>g>y>�>�>�>�>�>�>?"?8?T?f?x?�?�?�?�?�?   �   000=0^0t0�0�0�0�0�011G1t1�1�1"2*242F2P2k2�2�2�2�2�23=3f3�3�34'484A4T4�4�4�455*5<5b55�5�5d6y6�6�6�7�78!8D8d8�8�8�8�8949T9t9�9�9�9�9+:Q:�:;       _5A?a?�?�?     p   0E0�0�01R1�1�1�122e2�2�2%3b3�3�3�3"4U4�4�4%5u5�5�556u6�6%7�7�78U8�8�:�:>=�=�=�=�=�=�>�>�>�>b?p?�?�?   0 (  ^0l0�0�0�0�0�1
2#212�2�2�2�2�3�3�34434:4T4n4�4�4�4�4�4�4�4�4�45!5D5a5�5�5�56"6(6,62666<6@6F6J6O6U6Y6_6c6i6m6s6w6�6�6�6�6�6)7A7I7O7�7�7�7�788m8�899�9
:?:X:_:g:l:p:t:�:�:�:�:�:�:�:�:�: ;;N;T;X;\;`;�;�;�;�;�;�; <!<K<}<�<�<�<�<�<�<�<�<�<�<�<�<�<Q=[=h=�=�=�=w>�>�>�>�>�>??<?s?�?�?   @ �   M0_0�0�0�0�0�0h1�1�1�1�1`2r2�2�2�233!3,3�5S6�6�;�<D>�>�>�>�>�>�>�>????? ?'?.?5?<?C?J?R?Z?b?n?w?|?�?�?�?�?�?�?�?�?�?�?�?�?�?   P p  000/060J0Q0x0~0�0�0�0�0�0�0�0�0�0111 1,1:1@1L1R1_1i1p1�1�1�1�1�1�1	2I2O2y22�2�2�2S3v3�3�3�344"4.444D4J4_4m4x44�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4555555"515G5R5W5b5g5r5w5�5�5�5�5�5�5�56#6/6f6o6{6�6�6�6�6�6#7>7D7M7T7v7�7�7�7�7 888!8,858K8V8p8|8�8�8�8�8�8 9%90959S9�9�9�9	:*:0:b:�:�:;;3;L;�;�;�;!<'<K<i<�<�<�<�<�<7=B=L=]=h=?,?4?:???E?�?�?�?�?�?�? ` �   00F0�0�0�0�011(1-1a1f1t1|1�1�1�1�1�1�1�1�1�1�1�1
2�2�2�2�2q3�3�3�4�4�4�4K5e5�5�5�5�5�5�5�5�5�5�6�6�6�6�7�7�7�8�8�8959@9d9m9t9}9�9�9�9:4:G:_:q:�:�:=Q=�=a>q>}>�>�>�>�? p H   0�0,1x1�1�1�1�1H2p2u9�:�:%;�;�;�;-<q=�=�=�>�>�>?? ?�?�?�?�?   � �   00)050Z0c0l0y0�0�0�0�0�0�0�0�0�0111W1[1_1c1g1k1o1s1w1{11�1�1�1�1�12{2�2�2�2�2�2�2�23!3'303C3g3�34*4/4r6�6�6�6�6�6�6�6�6�6�677777<7B7M7R7Z7`7j7q7�7�7�7�7�7�7�7�7�7�7�7�7
8o8<<J<p<�<�<�>�>�>�>?3?F?{?�? � �   �0�011�1�2�2�233&3�3�34�5�5�5�5�5�5�5	6=6H6R6k6u6�6�6�67+7�7�7 8l8�8 99919L9T9\9s9�9�9�9�9�9�9�9�9$:5:X:;G;�;�;-<u<�<�<=?=n=�=R>\>i>�>�>�>?&? � �   ]0�031
2?2X2_2g2l2p2t2�2�2�2�2�2�2�2�2�2 33N3T3X3\3`3�3�3�3�3�3�3 4!4K4}4�4�4�4�4�4�4�4�4�4�4�4�4�4�7�9�9+:@:�:�:�:�: ;X;�;�;< <D<g<�<�<�<�<�=�=�=�=�=�=`>�>�>�>�>�>�>�>�>?S?X?�?�?�?�?�?�?   � h   )02080�0�0�0�01�1�1�233!31363N3T3c3i3x3~3�3�3�3�3�3�344;4�5�5�5�6�6
8�8�8�8P9c9~9�<�=C?r?�? � X   z1v3z3~3�3�3�3�3�3�3�4�6d88�8�8�89':�:�:-;{;�=�=�=�=�=�=!>N>`>m>y>�>�>�>�>�>�? � \   =0`0�0�172A2Y2`2j2r22�2�2O3�3�5�5�56)6;6M6_6q6�6�8�9�9`:B;�;�;�<�<�<9=P=�=�>�>�?   � H   �01%1�1�1�1}2�2�2Q3!686�9�9�9�9�9�9�9�9�9�9�9�9�9�:�:�:�:J;n;   � 4   x5 7�7�7	8#8,8�9�9�9�92:a:;;3<S<C=l=�=S?     �   30�0-1C1�1�1@2t2�2 3�3�3�3�3�3�3444&454A4N4r4�4�4�4�4�4
55"5F5u5�5�5�67U7r7�7�7�7�8�8R9Y=`=�=�=�=	>_>p>�>�>"?-?[?i?x?�?�?�?�?�?�?�?�?�?�?    `   0*0�0=1h1�1�1�1�1�1�1�2�2�23W3444!4(4:4�4C5o5�5�5�586u66�6�6�6#7�8�8�8�8�8�8�8�8     4   $1014181<1@1L1P1�4�4�4�4�4�5�5�6�6�6�6�6�7�7 0 �   �5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7 @ �   �2�2l3p3x3�3�3�3�3�3�3�3�3�3�3 444$44484H4L4T4l4|4�4�4�4�4�4�4�4585X5x5�5�5�5�5�5�566(6H6h6�6�6�6�67$7(7D7H7h7�7�7�7�7�7�78(8H8T8p8�8�8   P �   00P0T0X0\0`0d0h0l0�0�0�0�0�0�0�0�0�0�0�0�0 1111110141`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�142L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�344
444444"4&4*4.42464:4>4B4F4J4N4R4V4Z4^4b4f4j4n4r4v4z4~4�4�4�4X;P<�<�<�<�<�<=(=,=0=4=8=@=D=P=T=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?P?X?\?`?d?h?l?p?t?x?|?�?�?�? `    �2�2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        