MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       DT*� 5D� 5D� 5D��zҡ5D�	Mѡ5D�	Mǡt5D�'�?�5D� 5E�V5D�	M��A5D�	M֡5D�	Mա5D�Rich 5D�        PE  L <0N        � !	  N  �      �|     `                                                       � Y   �� (                            �    `a                            X� @            `                            .text   5M     N                   `.rdata  I1   `  2   R             @  @.data   X3   �     �             @  �.reloc  x)   �  *   �             @  B                                                                                                                                                                                                                                                                                                                                                                                                        U��E��dt���   uB��    ]á��H�Q4��+�=�  |� (  ���H�Q4�ң��   ]��������U����UV��H�AVR�Ѓ���^]� ��������������U���V��H�QV�ҡ��H�U�AVR�Ѓ���^]� U���V��H�QV�ҡ��U�H�E�IRj�PV�у���^]� ����������U����P�E�RP��VWP�EP�E�P�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ���������������U����P�R`��VW�E�P�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� �������U����H�U�I(��VWR�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]���U���8�EV�]�W�E3��]�3��E �]��3��U���  �E�E�M�E�P�M�Q�M��E�   �U��E�   �9  �U�R����<  ����u�E�PS�@C  ��������   V���=  �����   ���   jj���Ћ���tX�����   �E�Rlj P���҅�t;���D�ȋ��   ���$�ȋB0V�ЍM��(*  G���.���_�   ^��]ÍM��*  _3�^��]����U��QV�u���AM  �E���t}���$    ������   �ȋB��=/  t)-�  t"���=��t�����   �M��B(���'�����   �M��BL�ЍM�Q�.E  ������L  �E���u�^��]���������U��V�u��tB��I V�J��������   �B4������P����������   �B(�����Ћ���u�^]�U����H�A�� S�U�VR�Ћ��Q�J�E�P�ы��B�Pj j��M�h�aQ�ҍE�P�M�Q轊  �����B�P�M�Q���ҋu��$V��t@���H�Q�ҡ��H�Qj j�h�aV�ҡ��H�A�U�R�Ѓ���^[��]Ë��Q�B�Ћ��Q�J�E�VP�ы��B�P�M�Q�҃���^[��]��������������U���0  ���3ŉE�V�u���B�  ������Ph  � `��t������Q�������J�  �������jR誠  ��P����  ��������  �M���3�^�e ��]����U��Q����J  �E�����   ���$    ������   �ȋB�Ћ�=L  uN�Q@�E��J,P�у�h�  ���ի  ��u)�����   �M��PL�ҍE�P��B  �����ZJ  ������   �M��B(�ЉE����y�����]������U��V�u��t>��I �;��������   �B4����P����������   �B(�����Ћ���u�3�^]���諮  P����Y����U���`SV�uW����  �}�]��    ����  �����   �Bx���Ћ����   �E�Bx���Ћ��Q�M�RxQ���҅��w  �����   �B����=  ��   �����   �B����=  ��   ���QH�R`�E�P����� �]���@�]��@���PH�]��Rp�E�P��� �]Ћ��@�]��@���PH�]��Rh�E�P��� �]����@�]��@���]�h�  �E�W��E��X�E��X�;����EЃ����h�  �E�W�X�E��X�����E������h�  �E�W�X�E��X������� �����   �B4���ЋM�UWQRP�����   �B4����P�R��������   �B(�����Ћ����   ���B(���Ћ؅��=���_^[��]�������U��������   �SVW�}j j �������]������]��|�  P������]��;]�]�E���]�軴  �E�E���M��}���a�����]��$���  �M�Q��茿  �U�R��聿  j jjjj �����  �E�PVW����  P�����  P�U���C��;]�]~�����]�M���a�$�`�  �M�Q���%�  _��^[��]�������������U����P�B<��D�M�Ѕ�u���Q�J�EP�у�3���]Ë��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q���   ��j �E�Pj=�M�҅�u>���H�A�U�R�Ћ��Q�J�E�P�ы��B�P�MQ�҃�3���]ËM�V�E�PQj �U�R�M��������������Q�R�M�QP�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P<���M�ҋM�+�HPAQ�E�P�M�������Q�R�M�QP�ҡ��H�A�U�R�Ћ��Q�E�RP�M�Q�ҡ��H�A�U�R�Ћ��Qj j�h�a�E�P�J�ы��B�Px��(�M�Q�M��ҋ���H�A�ލU��RF�Ѓ���tB���Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�UR�Ѓ��   ^��]�j h�a�M���������Q�Rx�E�P�M��ҋ���H�A�ލU��RF�Ѓ���tB���Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�UR�Ѓ��   ^��]�j h�a�M��g������Q�Rx�E�P�M��ҋ���H�A�ލU��RF�Ѓ���tB���Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�UR�Ѓ��   ^��]�j h�a�M�������M�Q�M��V  �����B�P�M�Q�҃���tB���H�A�U�R�Ћ��Q�J�E�P�ы��B�P�MQ�҃��   ^��]�j h�a�M��j����E�P�M���  ���Q�J���E�P�ы��B�P�M܃�Q�ҡ��H�A�U�R�Ћ��Q�J�EP�у���t
�   ^��]�3�^��]�����������U���tSV3�W95�t)���jS���  ������uBF9<�����u܍M�l�  �M$�d�  ���B�P�M@Q�҃�_^�'  [��]Å�tˍEj P��  ����u1�M�%�  �M$��  ���Q�J�E@P�у�_^�'  [��]Ë��B�P�M�Q�ҡ��H�A3�Vj��U�h�aR�Ѓ��M�Q�M萇  �����B�P�M�Q�E��҃��}� �Mt-藄  �M$菄  ���H�A�U@R�Ѓ�_^�'  [��]�VjQ�u�賻  ���E��M;�u.�Q�  �M$�I�  ���B�P�M@Q�҃�_^�'  [��]ÍE�P�_�  �M�P覫  �M���  �M$覄  ����  �M$Q�M�"�  �M$�z�  Vh�a�M������U�R�M$耆  ���H�A�U�R�Ѓ��M$VQ蒑  ����t�U$VR���  ���M��v�  P�p����M����ŭ  �Mģ���  ���E�    ���   �R�E�Pj���ҋE����   ���Q@P�B,�Ћ�������   ���Q���   j j �E�P���ҡ��P�B0jh�  ���Ћ��Q�B0jh�  ���Ћ��Q�B0j h�  ���Ћ��Q�B0jh�  ���Ћ��Q�B0j h�  ���ЋEP�MT;�}Q�M�PQ��������E��U�j	R�l  �E�jP�tl  ���M�Q�M襃  Pj	�l  ���M��R�  ���B�P<�M@�҅�t"�E@P�M�豁  �M�Qj�Vl  ���M���  �E�Sj �U$RP��  ������t���Q���   j j V�M��ЍM�Qj	�l  �U�Rj�l  �E�P�ʸ  ���M�迁  �M�跁  �M���  �M见  �M$蟁  ���Q�J�E@P�у������_%����^'  [��]�Vh�a�M������M�Q�M$�)�  �����B�P�M�Q�E��҃��}� �x����M�,�  �M$�$�  ���H�A�U@R�Ѓ�_^�'  [��]�����U����  �  �E��E�P������ ���Q�������B�P<���M��҅���  ���H�A�U�R�Ћ��Q�Jj j��E�h�cP�эU�R�E�P�M�Q�a  �� P�M���  P�� ���R�����P���  ���M��V�  ���Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h�cP�эU�R�E�P�M�Q��  ��(P�M��i  P�� ���R������P�5�  ���M���  ���Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h�aP�ыE��='  ��  ��  ����  WPh�c��,�������j h�c������w���j h|c��<����e������:�EP�M�Q��e  ��P������WR�O�����P��,���P������Q�e  ����PR������P�!�����P�����Q��D���R�je  P��<���P������Q�  ��P��$���R�v  ��P������P�f  ��P��d���Q�V  ��P��4���R�F  ��P��T���P�6  ��P��t���Q�&  ��P������R�  ��P�M��
������H�A������R�Ћ��Q�J��t���P�ы��B�P��T���Q�ҡ��H�A��4���R�Ћ��Q�J��d���P�ы��B�P������Q�ҡ��H�A��$���R�Ћ��Q�J������P�ы��B�P��D���Q�ҡ��H�A������R�Ћ��Q�J������P�ы��B������Q�P�ҡ��H�A�U�R�Ћ��Q�J��<���P�ы��B�P�����Q�ҡ��H�A��,���R�Ѓ�@_��  j hTc�M��������Q�R�E�P�M�Q�ҡ��H�A�U�R�Ѓ��  �������0  �$��) j hc��\���������\���Q�M��F������B�P��\���Q�҃��A  j h�b��L����w�����L���P�M��������Q�J��L���P�у��  j h�b��l����9�����l���R�M���������H�A��l���R�Ѓ���   j h�b��|����������|���Q�M��������B�P��|���Q�҃��   j hTb�M�������E�P�M��U������Q�J�E�P�у��V���B�P�M�Q�ҡ��H�Aj j��U�h(bR�Ћ��Q�R�E�P�M�Q�ҡ��H�A�U�R�Ѓ� ���Q�J�E�P�ы��B�Pj j��M�h�aQ�ҡ��H�I�UR�E�P�ы��B�P�M�Q�ҡ��E�    �H���   h�ah�   h   �ҋ���,j �E��Qh   P�Bh�M���h1D4ChCD4Cjj j������Q�M��`  ���B�Pdj �M��ҋM�P�E�P�  �M��X  j�����Q������R�S�  ������j P�%�  �M�Q��  ���B�P�M�Q�҃���������y  �������y  �� �����y  ���H�A�U�R�ЍM�Q�~  ���E�    �B�P�MQ�҃���]��& 7' u' �' �' ��������U����   SVW�/~  h1D4ChCD4Cjj j�MQ�ȉE��Q~  ���B�P�M�Q�ҡ��H�Aj j��U�h�aR�Ћ��Q�J�E�P�ы��B�Pj j��M�h�aQ�ҡ��H�A��x���R�Ћ��Q�Jj j���x���h�aP�ы��B�P�M�Q�ҡ��H�A��@j j��U�h�aR�Ћ��Q�J�E�P�ы��B�Pj j��M�h�aQ�ҡ��E� �H�A�U�R�Ћ��Q�Jj j��E�h�aP�ы��B�P�M�Q�ҡ��H�Aj j��U�h�aR�ЋM���L3���}  ����  ����  3�3�j j�M�Q�M��+}  �E�<
�4  <�,  �M��}  ���� ;���  ;���  f�U����H�A��8���R�Ћ��Q�JV��8���jP�ы��B�P<���M��ҋ��Q�RLj�j���8���QP�M��ҡ��H�A��8���R�Ћ��B���M�Q�H����V�ы��B�P�M�VQ�҃���������wq�$�2 j h�a������
��������P�M��������Q�J�����P�у��/�U�R�M��!�M���M�Q��x�����U�R�M���M��E�P�R������Q�J��X���P�ы��B�Pj j���X���h�aQ�ҡ��H�I�U�R��X���P�ы��B�P��X���Q����  f�E����Q�J����(���P�ы��B�PV��(���jQ�ҡ��P�B<���M��Ћ��Q�RLj�j���(���QP�M��ҡ��H�A��(���R�Ѓ��j  ���B�M�Q�H����V�ы��B�P�M�VQ�҃�����������   �$�2 ���H�A��H���R�Ћ��Q�Jj j���H���h�aP�ы��B�@�M�Q��H���R�Ћ��Q�J��H���P�у� �h���B�@�M�Q�U�R���M�E��5���H�I��x���R�E�P���.���B�@�M�Q�U�R����E����Q�RP�M�Q�҃����H�A�U�R�Ћ��Q�Jj j��E�h�aP�ы��B�@�M�Q�U�R�Ћ��Q�J�E�P�у� �M�C�Ù�����z  ;��/���;��%����M��(y  �Uj R��  ���H�A��h���R�Ћ��Q�Jj j���h���h�aP�ы��B�P<���M��҅�uW���H�A�U�R�Ћ��Q�Jj j��E�h�cP�ы��B�@�M�Q�U�R�Ћ��Q�J�E�P�у� ���B�P<�M��҅�uW���H�A�U�R�Ћ��Q�Jj j��E�h�cP�ы��B�@�M�Q�U�R�Ћ��Q�J�E�P�у� ���B�PXj �M��ҋ���P�BXj �M��Ћ���h���QVP�B�H����V�ы��B�P��x���VQ�҃��E���P��q  ���U���R��q  ���������H�Q��D��V�ҡ��H�A��h���VR�Ѓ�W�2������Q�J��h���P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�E��JP�ы��B�P�M�Q�ҡ��H�A��x���R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҍE�P�uv  ��8�M�E�    �q  _^[��]ä, �, �, �, �, - :. �. �. �. �. �. ������������U���   SVW诵  �����p  ��I ���H�A�U�R�Ћ��Q�Jj j��E�h�cP�эU�R�;Y  ���H�A�U�R�Ћ��Q�J�E�P�ы��B�Pj j��M�h�cQ�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h�cP�у�D�U�R��`���P���\�  ���%q  ���Q�J���E�P�ы��B�@�M�Q�U�R�Ћ��Q���B<�M��Ћ��Qj�j�WP�BL�M��Ћ��Q�J�E�P�ы��B�@�M�Q�U�R�Ћ��Q�B<���M��Ћ��Q�RLj�j��M�QP�M��ҍE�P�X  ���Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�у���`����\o  ���B�P�M�Q�҃����p�  ���Q�J(P��|���P�ы����B�P�M�Q�ҡ��H�A�U�RW�Ћ��Q�J��|���P�эU�R�6W  ���H�A�U�R�Ћ����   �B(�� ���Ћ�����������Q�J�E�P�ы��B�Pj j��M�h�cQ�ҍE�P��V  ���Q�J�E�P�ы��B�P�M�Q�ҡ��H�Aj j��U�h�cR�ЍM�Q�V  ���B�P�M�Q�ҡ����   ���   ��j��jS藲  ��D����  �����   ���   ��3��Ѕ���  �����   ���   V���Ћ��Q�J���E�P�ы��B�Pj j��M�h�cQ�ҍE�P��U  ���Q�J�E�P�ы��B�P�M�Q�ҡ��H�Aj j��U�h�cR�Ћ��Q�J�E�P�ы��B�Pj j��M�h�cQ�҃�D��|���P��`���Q�����  ����m  ���E��B�P�M�Q�ҡ��H�U�R�I�E�P�ы��B�P<���M��ҋ��Q�M��RLj�j�QP�M��ҡ��H�A�U�R�Ћ��Q�R�E�P�M�Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҍE�P�T  ���Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J��|���P�у���`�����k  ���B�P�M�Q�҃�����  ���Q�J(P�E�P�ы����B�P�M�Q�ҡ��H�A�U�RW�Ћ��Q�J�E�P�эU�R��S  ���H�A�U�R�Ћ����   ���   �� ��F��;��w���_^[��]��������������U��E���   P������M�Q��������B�P<���M��҅�u"�M��k  ���H�A�U�R�Ѓ�3���]Ë��Q�J�E�P�ы��B�Pj j��M�h dQ�ҍE�P�M�Q�U�R�  �� P��|����j  P�E�P�M�Q��m  ����|����j  ���B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�Pj j��M�h�cQ�҃��E�P�M���j  P�M�Q�U�R��   P�_R  ���H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҍE�j P�w  ��$��tZ���B�P�M�Q�ҡ��H�Aj j��U�h�cR�ЍM�Q��Q  ���B�P�M�Q�ҍE���P�6i  �������M��fi  �M��^i  ���Q�J�E�P�у�3���]����U����P�E�RxP�����@]� ���U����H�QV�uV�ҡ��H�U�AVR�Ћ��Q�B<�����Ћ��Q�M�RLj�j�QP���ҋ�^]��������̡��  �����  ;��@����������U������ ��������  v3���]Ë@�P�M�Q�ҡ��H�Aj j��U�hLdR�ЍM�Q�P  ���B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�Jj j��E�hdP�эU�R�YP  ���H�A�U�R�Ѓ�8�   ��]�����������������������������U����  ���=�  v3�]ËE�� t��t-Vu�u��]����   ]ù ��ܿ  �����]�����U��E��� ]��h�PhD �0�  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h�jhD �\�  ����t
�@��t]��3�]��������Vh�j\hD ���,�  ����t�@\��tV�Ѓ���^�����Vh�j`hD �����  ����t�@`��tV�Ѓ�^�������U��Vh�jdhD �����  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�jhhD ����  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�jlhD ���L�  ����t�@l��tV�Ѓ�^�������U��Vh�h�   hD ����  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h�   hD �����  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�jphD ���y�  ����t�@p��t�MQV�Ѓ�^]� ��^]� ��U��Vh�jxhD ���9�  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�jxhD �����  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�jxhD ����  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������h�jhD �_�  ����t	�@��t��3��������������U��V�u�> t+h�jhD �#�  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h�jhD ���  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�jhD ����  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�jhD ���Y�  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�j hD ����  ����t�@ ��tV�Ѓ�^�3�^���Vh�j$hD ����  ����t�@$��tV�Ѓ�^�3�^���U��Vh�j(hD ��蹿  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�j,hD ���i�  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�j(hD ���)�  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�j4hD ���ܾ  ����t�@4��tV�Ѓ�^�3�^���U��Vh�j8hD ��詾  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�j<hD ���Y�  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�jDhD ����  ����t�@D��tV�Ѓ�^�3�^���U��Vh�jHhD ����  ����t�M�PHQV�҃�^]� U��Vh�jLhD ��蹽  ����u^]� �M�PLQV�҃�^]� �����������U��Vh�jPhD ���y�  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�jThD ���<�  ����u^Ë@TV�Ѓ�^���������U��Vh�jXhD ���	�  ����t�M�PXQV�҃�^]� U��Vh�h�   hD ���ּ  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�h�   hD ��膼  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�h�   hD ���6�  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD �����  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ��趻  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���v�  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�h�   hD �5�  ����u���H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]��U��Vh�h�   hD ��覺  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�h�   hD ���V�  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   hD ����  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   hD ���ֹ  ����t���   ��t�MQ����^]� 3�^]� �Vh�h�   hD ��虹  ����t���   ��t��^��3�^����������������U��Vh�h�   hD ���V�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�h�   hD ����  ����t���   ��t�MQ����^]� ��������U��Vh�h�   hD ���Ƹ  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh�h�   hD ���y�  ����t���   ��t��^��3�^����������������VW��3����$    �h�jphD �/�  ����t�@p��t	VW�Ѓ�����8 tF��_��^�������U��SW��3�V��    h�jphD �߷  ����t�@p��t	WS�Ѓ�����8 tqh�jphD 護  ����t�@p��t�MWQ�Ѓ������h�jphD �{�  ����t�@p��t	WS�Ѓ����V���7�����tG�]����E^��t�8��~=h�jphD �.�  ����t�@p��t	WS�Ѓ�����8 u_�   []� _3�[]� ����������U��Vh�j\hD ���ٶ  ����t3�@\��t,V��h�jxhD 跶  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�j\hD ���y�  ����t3�@\��t,V��h�jdhD �W�  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�j\hD ����  ����tG�@\��t@V�ЋEh�jdhD �E��E�    �E�    ��  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�j\hD ��虵  ����t\�@\��tUV��h�jdhD �w�  ����t�@d��t
�MQV�Ѓ�h�jhhD �N�  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�j\hD ���	�  ������   �@\��t~V��h�jdhD ��  ����t�@d��t
�MQV�Ѓ�h�jhhD 躴  ����t�@h��t
�URV�Ѓ�h�jhhD 葴  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�jthD ���V�  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�j`hD ��  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh����_�����^��]� ������U���Vh�h�   hD ���ó  ����tR���   ��tH�MQ�U�R���ЋuP������h�j`hD 芳  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t�����   P�B@��]� �E��t�����   P�BD��]� �����   R�PD��]� �����U����P@�Rd]�����������������U����P@�Rh]�����������������U����P@�Rl]�����������������U����P@�Rp]�����������������U������   ���   ]�����������U������   ���   ]����������̡��P@�Bt����̡��P@�Bx�����U����P@�R|]����������������̡��P@���   ������   �Bt��U����P@���   ]�������������̡��P@���   ��U����P@���   ]��������������U����P@���   ]��������������U����P@���   ]��������������U����P@���   ]��������������U���V��H@�QV�ҋM����t��#������Q@P�BV�Ѓ�^]� �̡��PH���   Q�Ѓ�������������U����P@�EPQ�JL�у�]� ���̡��P@�BHQ�Ѓ����������������U����P@�EP�EP�EPQ�J�у�]� ������������U����P@�EPQ�J�у�]� ����U����P@�EP�EPQ�J�у�]� U����P@�EPQ�J �у�]� ����U������   �R]��������������U������   �R]��������������U������   �R ]��������������U������   ���   ]�����������U������   ��D  ]�����������U����E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U������   ���   ]����������̡����   �B$����H@�Q0�����U����H@�A4j�URj �Ѓ�]����U����H@�A4j�URh   @�Ѓ�]�U����H@�U�E�I4RPj �у�]�̡��H|�������U��V�u���t���Q|P�B�Ѓ��    ^]��������̡��H|�Q �����U��V�u���t���Q|P�B(�Ѓ��    ^]��������̡��H@�Q0�����U��V�u���t���Q@P�B�Ѓ��    ^]���������U����H@���   ]��������������U��V�u���t���Q@P�B�Ѓ��    ^]��������̡��PH���   Q�Ѓ�������������U����PH�EPQ��d  �у�]� �U����H �IH]�����������������U��}qF uHV�u��t?�����   �BDW�}W���Ћ��Q@�B,W�Ћ��Q�M�Rp��VQ����_^]����������̡��P@�BT�����U����P@�RX]�����������������U����P@�R\]����������������̡��P@�B`�����U����H��T  ]��������������U����H@�U�A,SVWR�Ћ��Q@�J,���EP�ы��Z��h��hE  �΋��l  Ph��hE  ���l  P��T  �Ѓ�_^[]����U������   ���   ]�����������U����H@�AV�u�R�Ѓ��    ^]��������������U����PL�E��  PQ�MQ�҃�]� ������������̡��PD�BQ�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�BQ�Ѓ����������������U����PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U����PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U����PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U����PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U����PX�EPQ�J�у�]� ����U����PX�EPQ�J�у�]� ����U����PX�EPQ�J�у�]� ����U����PX�EPQ�J�у�]� ����U����PX�EPQ�J$�у�]� ����U����PX�EPQ�J �у�]� ����U����PD�EP�EPQ�J�у�]� U����HD�U�j R�Ѓ�]�������U����H@�AV�u�R�Ѓ��    ^]��������������U����HD�	]��U����H@�AV�u�R�Ѓ��    ^]��������������U����HD�U�j R�Ѓ�]�������U����H@�AV�u�R�Ѓ��    ^]��������������U����U�HD�Rh'  �Ѓ�]����U����H@�AV�u�R�Ѓ��    ^]�������������̡��HD�j h�  �҃�����������U����H@�AV�u�R�Ѓ��    ^]�������������̡��HD�j h:  �҃�����������U����H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E������   �R�E�Pj�����#E���]�̡��HD�j h�F �҃�����������U����H@�AV�u�R�Ѓ��    ^]�������������̡��HD�j h�_ �҃�����������U����H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E����E�    ���   �R�E�Pj������؋�]� ̡��PD�B$Q�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ����������������U����E�PH�B���$Q�Ѓ�]� ���������������U����PH�EPQ���   �у�]� �U����PH�EPQ���  �у�]� �U����PH�EPQ���  �у�]� �U����PH�EP�EPQ��  �у�]� �������������U����PH�EP�EPQ��  �у�]� ������������̡��PH���  Q�Ѓ�������������U����PH�EPQ���  �у�]� ̡��PH���   j Q�Ѓ�����������U����PH�EPj Q���   �у�]� ��������������̡��PH���   jQ�Ѓ�����������U����PH�EPjQ���   �у�]� ��������������̡��PH���   jQ�Ѓ����������U����PH�EPjQ���   �у�]� ���������������U����PH�EP�EPQ���   �у�]� �������������U����PH�EP�EPQ���   �у�]� ������������̡��PH���   Q�Ѓ�������������U����PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP�������������t�E���QH���   PVW�у���_^]� �����U��EVW���MPQ�����������t�M���BH���   QVW�҃���_^]� ̡��PH���   Q�Ѓ������������̡��PH���   Q�Ѓ�������������U����PH�EPQ���   �у�]� �U����PH�EPQ���   �у�]� �U����PH�EP�EPQ��8  �у�]� �������������U����PH�EP�EPQ��   �у�]� ������������̡��PH���  Q�Ѓ������������̡��PH���  Q�Ѓ������������̡��PH���  Q�Ѓ������������̡��PH��  Q�Ѓ������������̡��PH��  Q�Ѓ�������������U����PH�EP�EPQ��  �у�]� �������������U����PH�EP�EP�EPQ��   �у�]� ���������U����PH�EP�EP�EP�EPQ��|  �у�]� �����U����PH�EPQ��  �у�]� ̡��PH��T  Q�Ѓ�������������U����PH�EP�EPQ��  �у�]� �������������U����PH�EPQ��8  �у�]� �U����PH�EPQ��<  �у�]� �U����PH�EPQ��@  �у�]� �U����PH�EP�EP�EPQ��D  �у�]� ��������̡��PH��L  Q��Y��������������U����PH�EPQ��H  �у�]� ̡�V��H@�Q,WV�ҋ��Q��j �ȋ��   h�  �Ћ��QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡��P@�B,Q�Ћ��Q��j �ȋ��   h�  �������U����E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U����E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U����PH�EP�EP�EPQ��   �у�]� ��������̡��HH��  ��U����HH��  ]��������������U����E�PH��$  ���$Q�Ѓ�]� �����������̡��PH��(  Q�Ѓ�������������U����PH�EP�EPQ��,  �у�]� �������������U����E�PH�EP�E���$PQ��0  �у�]� ���̡��PH���  Q�Ѓ������������̡��PH��4  Q�Ѓ������������̋��     �������̡��PH���|  jP�у���������U����UV��HH��x  R��3Ƀ������^��]� ��̡��PH���|  j P�у��������̡��PH��P  Q�Ѓ������������̡��PH��T  Q�Ѓ������������̡��PH��X  Q�Ѓ�������������U����PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡��PH��`  Q�Ѓ�������������U����PH�EPQ��d  �у�]� �U����E�PH��h  ���$Q�Ѓ�]� ������������U����E�PH��t  ���$Q�Ѓ�]� ������������U����E�PH��l  ���$Q�Ѓ�]� ������������U����PH�EPQ��p  �у�]� �U����PH�EP�EP�EP�EPQ���  �у�]� �����U����PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U����E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E���HH�E���   R�U���$P�ERP�у�]����������������U���E�M��d� �M;�|�M;�~��]�����������U����PH�E���   Q�MPQ�҃�]� ������������̡��PH���   Q��Y�������������̡��PH���   Q�Ѓ������������̡��PH���   Q��Y��������������U����PH�EP�EPQ���   �у�]� �������������U����PH�EP�EP�EP�EP�EPQ���  �у�]� ̡��PH��t  Q��Y�������������̋�� �d�@    ���d���Pl�A�JP��Y��������U���V��Hl�V�AR�ЋE����u
�   ^]� ���Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË��QlP�B�Ѓ�������U����Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E���HH�ER�U���$P���  R�Ѓ�]����U����HH���  ]��������������U����HH���  ]��������������U��U0�E(���HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U����HH���  ]��������������U����E�PH�EP���$Q���  �у�]� ��������U���SV����  �؉]����   �} ��   ���HH��p  j h�  V�҃��E��u
^��[��]� �MW3��}���  ����   �]��I �E�P�M�Q�MW诔  ��ta�u�;u�Y�I ������u�E�������L�;Ht-���Bl�S�@����QR�ЋD������t	�M�P蓓  F;u�~��}��MG�}��^�  ;��v����]�_^��[��]� ^3�[��]� ��������������U�����SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u���HH���  �'��u���HH���  ���uš��HH���  S�ҋȃ��E��t�W�$�  ���HH���   h�  S3��҃����  ���_�u����    ���Hl�U�B�IWP�ы�������   ���F�J\�UP�A,R�Ѓ���t�K�Q�M�E�  ���F�J\�UP�A,R�Ѓ���t�K�Q�M��  �E��;Pt&�F���Q\�J,P�EP�у���t	�MS��  ���v�B\�M�P,VQ�҃���t�M�CP�Ñ  ���QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U����HH���   ]�������������̡��PH���   Q��Y��������������U����HH���  ]��������������U�����P���   V�uW�}���$V�����E������At���E������z����؋��Q�B,���$V����_^]����������������U���0����U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١��]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U����HH�]��U����H@�AV�u�R�Ѓ��    ^]�������������̡��HH�h�  �҃�������������U����H@�AV�u�R�Ѓ��    ^]��������������U����HH�Vh  �ҋ�������   �EPh�  � �������t]���QHj P���   V�ЋMQh(  ���������t3���JH���   j PV�ҡ����   �B��j j���Ћ�^]á��H@�QV�҃�3�^]�������U����H@�AV�u�R�Ѓ��    ^]��������������U����HH�Vh�  �ҋ�����u^]á��HH�U�E��  RPV�у���u���B@�HV�у�3���^]�������U����H@�AV�u�R�Ѓ��    ^]��������������U����HH�I]�����������������U����H@�AV�u�R�Ѓ��    ^]��������������U����PH�EPQ���  �у�]� �U����PH�EPQ���  �у�]� ̡��PH���  Q�Ѓ�������������U����HH���  ]��������������U����E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡��PH���  Q�Ѓ�������������U����PH�EP�EPQ���  �у�]� ������������̡��PH��  Q�Ѓ�������������U����PH�EP�EP�EPQ���  �у�]� ��������̡��PH���  Q�Ѓ������������̡��PH���  Q�Ѓ�������������U����PH�EPQ��  �у�]� �U����PH�EPQ��  �у�]� ̋������������������������������̡��HH���  ��U����HH���  ]��������������U����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡��PH��,  Q�Ѓ�������������U����PH�EPQ��X  �у�]� ̡��PH��\  Q�Ѓ�������������U����HH��0  ]��������������U�����W���HH���   j h�  W�҃��} u�   _��]� Vh�  ������������   ���HH���   j VW�҃��M��H  ���P�E�R0Ph�  �M����E���P�B,���$h�  �M��Ћ��Q@�J(j �E�PV�у��M��H  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7���U�HH���   RW�Ѓ���u���QH���   jW�Ѓ���t�   �����   ���QH���   W�Ѓ��} u(���E�QH�M���  P�ESQ�MPQW�҃��B�u��t;���U�HH�ER�USP���  VRW�Ћ����   �B(�����Ћ���uŃ; u���QH���   W�Ѓ���t3���   �W��u1���QH���   �Ћ��E�QH���   PW�у�_^[]� ���BH���   �у��} u0���M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ���QH�h  �Ћ؃���u_^[]� �����   �u�Bx���Ћ����   P�B|���Ѕ�tU���E�QH�MP�Ej Q���  VPW�у���t�����   �ȋBHS�Ћ����   �B(���Ћ���u�_^��[]� ��������������U��EV���u���HH���  �'��u���HH���  ���u���HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D���HH���   S�]VWh�  S�ҋ���HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��.
  �����   �B���Ћ�=�  ��  �QH���   Wh:  S�Ћ��QH�E����   h�  S�Ћ��QHW�����   h�  S�uԉ}��Ћ��QH�E苂  S�Ћ��QH�EЋ��  S�Ѓ�(�E��E��d��~~�M���M�I �MЅ�tMj�W�1�  ���t@�@�Ẽ|� �4�~����%�������;�u/���@�  ;E�~�E؋���  E���E�;Pu�E���E��E�G;}�|��}� tv�u�j S����������  ���������tV���1����}�;�uK���H���  �4�h�d��h�  V�҃��E���N  �M�PVP����P�  ����}ܡ��H���  �4�h�d��h�  V�҃��E����  �M�3�;�t;�tVQP�H  ���E�;�~-���Qh�d��h�  P���   �Ѓ��E�;���  ���E��QH��  j�PS�у�����  �u�;�tjS���}������{  ��������E���}���BH���   Wh�  S�у�3�9}ԉE�}��`  �}���}Ȑ�MЅ��R  �U�j�R�:�  ����>  �M̍@�|� ���]�~����%�������9E���  ����  �E�3�3�9C�E܉M���   ��$    �����������tk�]��}������������ϋ9�<��}�@�҉��y�]��|��]�@@�z�<��y�]��|��]�@@�z�<��I�}��]�@���M��}�@����@�M�A;K�M��t����E؅��9  �+U�j��PR�M�襉  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$�� �U����4�"�M����t��U����t�
�M����t�M���;]�|��E܃�F;]؉M��	����U�;U��
  �U�R��g  �E�P��g  �M�Q��g  ��_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���P�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@��;EԉE��}�������U�R��e  �E�P�e  ���  ���   �B����=  ��  ���QH���   j h(  S�Ћ��QH�����   h(  S�ЋЃ�3��U؅�~'����    �ǅ�t�|� t�4N��tN�@;�|�u��u܋��Q���  �4v�h�d��hK  V�Ѓ��E�����   �M��t��tVQP�X�  ���u؋��Q���  �h�d��hP  V�Ѓ��E���tP��t��tVWP��  ���M����+��RH��PQ�E���   S�Ѓ���u�M�Q�rd  �U�R�id  ��_^3�[��]á��HH���   j h�  S�҉E����HH���   j h(  S��3�3���3�9]؉E��}ĉ]��7  �U��څ��  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�F@F����;�|��}ă|� ts�U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�F�v�Ћ��A�B�A�B�A�B�A�B�I�J�U�F<ډ}�C;]؉]�������M�3�3�;�~�U����$    ��t���   @;�|��U�R�b  ���E�P�b  ��_^�   [��]�_� j� v� �� ������������U��U��t�M��t�E��tPRQ���  ��]������������U��E� �M+]� ���������������U��V��V��d���Hl�AR�Ѓ��Et	V�4e  ����^]� ����������U����P8�EPQ�JD�у�]� ���̡��H8�Q<�����U����H8�A@V�u�R�Ѓ��    ^]�������������̡��H8�������U����H8�AV�u�R�Ѓ��    ^]��������������U����P8�EP�EP�EPQ�J�у�]� ������������U����P8�EP�EPQ�J�у�]� ���P8�BQ�Ѓ����������������U����P8�EPQ�J �у�]� ����U����P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U����P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U����P8�EP�EPQ�J(�у�]� U����P8�EP�EP�EPQ�J,�у�]� ������������U����P8�EP�EP�EPQ�J�у�]� ������������U����P8�EP�EP�EP�EP�EPQ�J�у�]� ����U����P8�EP�EPQ�J0�у�]� U����P8�EP�EP�EPQ�J4�у�]� ������������U����P8�EPQ�J8�у�]� ����U����H��x  ]��������������U����H��|  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H�A,]�����������������U����H�QV�uV�ҡ��H�Q8V�҃���^]�����̡��H�Q<�����U����H�I@]����������������̡��H�QD����̡��H�QH�����U����H�AL]�����������������U����H�IP]�����������������U����H��<  ]��������������U����H��,  ]��������������U����H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡��H���   ����H���  ��U����H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U����H�A]�����������������U����H��\  ]��������������U����H�AT]�����������������U����H�AX]�����������������U����H�A\]����������������̡��H�Q`����̡��H�Qd����̡��H�Qh�����U����H�Al]�����������������U����H�Ap]�����������������U����H�At]�����������������U����H��D  ]��������������U����H��  ]��������������U����H�Ix]�����������������U����H��@  ]��������������U��V�u���  ���H�U�A|VR�Ѓ���^]���������U����H���   ]��������������U����H��h  ]��������������U����H��d  ]��������������U����H���  ]�������������̡��H���   ��U����H��l  ]��������������U����H��   ]��������������U����H��  ]��������������U��V�u���B2  ���H���   V�҃���^]���������̡��H��`  ��U����H��  ]��������������U����H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U����H���  ]��������������U��U�E���H�E���   R���\$�E�$P�у�]�U����H���   ]��������������U����H���   ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���   ]��������������U����H���   ]��������������U����H���   ]��������������U����H���   ]��������������U����H���   ]��������������U����H���   ]��������������U����P���E�P�E�P�E�PQ���   �у����#E���]����������������U����P���E�P�E�P�E�PQ���   �у����#E���]����������������U����P���E�P�E�P�E�PQ���   �у����#E���]����������������U����H��8  ]��������������U��V�u(V�u$�E�@���R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@���R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U����P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U����P0�EP�EP�EP�EPQ���   �у�]� ����̡��P0���   Q�Ѓ�������������U����P0�EP�EPQ���   �у�]� �������������U����P0�EP�EP�EP�EPQ���   �у�]� ����̡��P0���   Q�Ѓ������������̡��H0���   ��U����H0���   V�u�R�Ѓ��    ^]�����������U����H��H  ]��������������U����H��T  ]�������������̡��H��p  ����H���  ��U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �����   �Qj PV�ҡ����   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M��+  P�E�hicMCP�k������M���+  �����   �JT�E�P�у���u(�u���Z+  �����   ��M�Q�҃���^��]á����   �AT�U�R�Ћu��P���Z+  �����   �
�E�P�у���^��]�������������U����H��  ]��������������U����H��\  ]��������������U����H�U��t  ��V�uVR�E�P�у�����  �M��  ��^��]�����U����H�U���  ��VWR�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]����������������U����H�U���  ��VWR�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]����������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H�U�E��VWj R�UP�ERP��t  �U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�(_��^��]��U����H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �����   j P�BV�Ћ����   �
�E�P�у�$��^��]���U����H��8  ]��������������U���  ���3ŉE��M�EPQ������h   R�� ����|	=�  |#����H��0  h�dhF  �҃��E� ���H��4  ������Rh,e�ЋM�3̓��>�  ��]�������U����H��  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]����U����H��  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]����U����H��p  ��$�҅�trh���M��&  ���P�E�R4Ph���M��ҡ��P�E�R4Ph���M���j �E�P�M�hicMCQ���������   ��M�Q�҃��M��t&  ��]�U����H��p  ��$V�҅�u���H�u�QV�҃���^��]�Wh!���M���%  ���P�E�R4Ph!���M���j �E�P�M�hicMCQ���������   �QHP�ҋu�����H�QV�ҡ��H�QVW�ҡ����   ��U�R�Ѓ�$�M��%  _��^��]������U����H��p  ��$V�҅�u���H�u�QV�҃���^��]�Wh����M��%  ���P�E�R4Ph����M���j �E�P�M�hicMCQ���������   �QHP�ҋu�����H�QV�ҡ��H�QVW�ҡ����   ��U�R�Ѓ�$�M���$  _��^��]������U����H��p  ��$�҅�u��]�Vh#���M��d$  ���P�E�R4Ph#���M���j �E�P�M�hicMCQ����������   �Q8P�ҋ�����   ��U�R�Ѓ��M��E$  ��^��]���������������U����H��p  ��$�҅�u��]�Vhs���M���#  ���P�E�R4Phs���M���j �E�P�M�hicMCQ�W��������   �Q8P�ҋ�����   ��U�R�Ѓ��M��#  ��^��]���������������U����H���  ]��������������U����H��@  ]��������������U����H���  ]��������������U��V�u���t���QP��D  �Ѓ��    ^]������U����H��H  ]��������������U����H��L  ]��������������U����H��P  ]��������������U����H��T  ]��������������U����H��X  ]��������������U����H��\  ]�������������̡��H��d  ��U����H��h  ]��������������U����H��l  ]�������������̡��H���  ��U����H�U���  ��VR�E�P�ыu��P���!  �M��!  ��^��]�����U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H��$  ]��������������U����H��(  ]��������������U����H��,  ]�������������̡��H��0  ����H��<  ��U����H���  ]�������������̡��H���  ��U����H���  ]������������������������������U����H��  ]�������������̡��H��P  ������   ���   ��Q��Y��������U����H�A�U��� R�Ћ��Q�Jj j��E�h0eP�ыUR�E�P�M�Q�=������B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�у�,��]��U����P�EP�EP�EPQ�J�у�]� �����������̡�V��H�QV�ҡ��H$�QDV�҃���^�����������U���V��H�QV�ҡ��H$�QDV�ҡ��U�H$�AdRV�Ѓ���^]� ��U���V��H�QV�ҡ��H$�QDV�ҡ��U�H$�ARV�Ѓ���^]� ��U���V��H�QV�ҡ��H$�QDV�ҡ��H$�U�ALVR�Ѓ���^]� �̡�V��H$�QHV�ҡ��H�QV�҃�^�������������U����P$�EPQ�JL�у�]� ����U����P$�R]�����������������U����P$�Rl]����������������̡��P$�Bp����̡��P$�BQ�Ѓ����������������U����P$��VWQ�J�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]� ���U����P$�EPQ�J�у�]� ����U����P$��VWQ�J �E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]� ���U����P$��VWQ�J$�E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e������Q$�JH�E�P�ы��B�P�M�Q�҃���^��]� ����̡��P$�B(Q��Yá��P$�BhQ��Y�U����P$�EPQ�J,�у�]� ����U����P$�EPQ�J0�у�]� ����U����P$�EPQ�J4�у�]� ����U����P$�EPQ�J8�у�]� ����U����UV��H$�ALVR�Ѓ���^]� ��������������U����H�QV�uV�ҡ��H$�QDV�ҡ��H$�U�ALVR�Ћ��E�Q$�J@PV�у���^]�U����UV��H$�A@RV�Ѓ���^]� ��������������U����P$�EPQ�J<�у�]� ����U����P$�EPQ�J<�у����@]� ���������������U����P$�EP�EPQ�JP�у�]� U����P$�EPQ�JT�у�]� ���̡��H$�QX�����U����H$�A\]�����������������U����P$�EP�EP�EPQ�J`�у�]� �����������̡��H(�������U����H(�AV�u�R�Ѓ��    ^]��������������U����P(�R]����������������̡��P(�B�����U����P(�R]�����������������U����P(�R]�����������������U����P(�R ]�����������������U����P(�E�RjP�EP��]� ��U����P(�E�R$P�EP�EP��]� ���P(�B(����̡��P(�B,����̡��P(�B0�����U����P(�R4]�����������������U����P(�RX]�����������������U����P(�R\]�����������������U����P(�R`]�����������������U����P(�Rd]�����������������U����P(�Rh]�����������������U����P(�Rx]�����������������U����P(�Rl]�����������������U����P(�Rt]�����������������U����P(�Rp]�����������������U������E�    �E�    �P(�RhV�E�P���҅���   �E���uG���H�A�U�R�Ћ��Q�E�RP�M�Q�ҡ��H�A�U�R�Ѓ��   ^��]� ���Qh4eh8  P���   �Ћ����E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P��<  ��3�^��]� �M��U�j IQ�MR�����E�P��<  ���   ^��]� ���������������U�����V��H�A�U�R�Ѓ��M�Q������^��u���B�P�M�Q�҃�3���]� ���H$�E�I�U�RP�ы��B�P�M�Q�҃��   ��]� �U��Q���P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U����P(�R8]�����������������U����P(�R<]�����������������U����P(�R@]�����������������U����P(�RD]�����������������U����P(�RH]�����������������U����P(�E�R|P�EP��]� ����U����P(�RL]�����������������U����E�P(�BT���$��]� ���U����E�P(�BPQ�$��]� ����̡��H(�Q�����U����H(�AV�u�R�Ѓ��    ^]��������������U����P(���   ]��������������U����H(�A]����������������̡��H,�Q,����̡��P,�B4�����U����H,�A0V�u�R�Ѓ��    ^]�������������̡��P,�B8�����U����P,�R<��VW�E�P�ҋu�����H�QV�ҡ��H$�QDV�ҡ��H$�QLVW�ҡ��H$�AH�U�R�Ћ��Q�J�E�P�у�_��^��]� �������U����P,�E�R@��VWP�E�P�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ��̡��H,�j j �҃��������������U����P,�EP�EPQ�J�у�]� U����H,�AV�u�R�Ѓ��    ^]�������������̡��P,�B����̡��P,�B����̡��P,�B����̡��P,�B ����̡��P,�B$����̡��P,�B(�����U����P,�R]�����������������U����P,�R��VW�E�P�ҋu�����H�QV�ҡ��H$�QDV�ҡ��H$�QLVW�ҡ��H$�AH�U�R�Ћ��Q�J�E�P�у�_��^��]� �������U����H��D  ]��������������U����H��H  ]��������������U����H��L  ]��������������U����H�I]�����������������U����H�A]�����������������U����H�I]�����������������U����H�A]�����������������U����H�I]�����������������U����H���  ]��������������U����H�A]�����������������U���V�u�E�P���k������Q$�J�E�P�у���u-���B$�PH�M�Q�ҡ��H�A�U�R�Ѓ�3�^��]Ë��Q�J�E�jP�у���u=�U�R��������u-���H$�AH�U�R�Ћ��Q�J�E�P�у�3�^��]Ë��B�HjV�у���u���B�HV�у����I������Q$�JH�E�P�ы��B�P�M�Q�҃��   ^��]�����������U����H�A ]�����������������U����H�I(]�����������������U����H��  ]��������������U����H��   ]��������������U����H��  ]��������������U����H��  ]��������������U����H�A$��V�U�WR�Ћ��Q�u���BV�Ћ��Q$�BDV�Ћ��Q$�BLVW�Ћ��Q$�JH�E�P�ы��B�P�M�Q�҃�_��^��]������U����H���  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q$�BDV�Ћ��Q$�BLVW�Ћ��Q$�JH�E�P�ы��B�P�M�Q�҃�_��^��]���U����H���  ]��������������U���<��SVW�E�    ��t�E�P�   �X������/���Q�J�E�P�   �ы��B$�PD�M�Q�҃��}���H�u�QV�ҡ��H$�QDV�ҡ��H$�QLVW�҃���t)���H$�AH�U�R����Ћ��Q�J�E�P�у���t&���B$�PH�M�Q�ҡ��H�A�U�R�Ѓ�_��^[��]���U����H�U���  ��VWR�E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡��H���   ��U����H���   V�uV�҃��    ^]�������������U����P�]����P�B����̡��P���   ��U����P�R`]�����������������U����P�Rd]�����������������U����P�Rh]�����������������U����P�Rl]�����������������U����P�Rp]�����������������U����P�Rt]�����������������U����P���   ]��������������U����P�Rx]�����������������U����P���   ]��������������U����P�R|]�����������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P�EPQ��  �у�]� �U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U��E��t ���R P�B$Q�Ѓ���t	�   ]� 3�]� U����P �E�RLQ�MPQ�҃�]� U��E��u]� ���R P�B(Q�Ѓ��   ]� ������U����P�R]�����������������U����P�R]�����������������U����P�R]�����������������U����P�R]�����������������U����P�R]�����������������U����P�R]�����������������U����P�E�R\P�EP��]� ����U����E�P�B ���$��]� ���U����E�P�B$Q�$��]� �����U����E�P�B(���$��]� ���U����P�R,]�����������������U����P�R0]�����������������U����P�R4]�����������������U����P�R8]�����������������U����P�R<]�����������������U����P�R@]�����������������U����P�RD]�����������������U����P�RH]�����������������U����P�RL]�����������������U����P�RP]�����������������U����P���   ]��������������U����P�RT]�����������������U����P�EPQ��  �у�]� �U����P���   ]��������������U����P���   ]��������������U����P�RX]����������������̡��P���   ��U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]�������������̡��P���   ��U����P���   ]�������������̡��P���   ����P���   ����P���   ��U����H���   ]��������������U����H��   ]��������������U����H�U�E��VWRP���  �U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]������������U����H���  ]��������������U����P(�} �R8����P��]� �U����P�BdS�]VW��j ���Ћ��Q�����   h4eFhc  V�Ћ����E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ��Q(�BHV���Ѕ�t ���Q(�E�R VP���҅�t�   �3��EP�(  ��_��^[]� ������U���V�E���MP�{���P���#������Q�J���E�P�у���^��]� ��̡��P�BVj j����Ћ�^���������U����P�E�RVj P���ҋ�^]� U����P�E�RVPj����ҋ�^]� ���P�B�����U����P���   Vj ��Mj V�Ћ�^]� �����������U����P�EPQ�J�у�]� ����U����P�EPQ�J�у����@]� ���������������U����P�E�RtP�ҋ����   P�BX�Ѓ�]� ���U����P�E�Rlh#  P�EP��]� ���������������U����P�E�RlhF  P�EP��]� ���������������U����P�E�RtP�ҋ����   �M�R`QP�҃�]� ���������������U����P���   ]��������������U����P�E���   P�҅�u]� �����   P�B�Ѓ�]� �������̡��HL���   ��U����H@�AV�u�R�Ѓ��    ^]�������������̡��HL�������U����H@�AV�u�R�Ѓ��    ^]�������������̡��PL���   Q�Ѓ�������������U����PL�EP�EPQ���   �у�]� �������������U���V��HL���   V�҃���u���U�HL���   j RV�Ѓ�^]� �����   �ȋBP�Ћ����   �MP�BH��^]� �����̡��PL��(  Q�Ѓ�������������U����PL�EP�EPQ��,  �у�]� ������������̡��HL�Q�����U����H@�AV�u�R�Ѓ��    ^]��������������U����PL�E�R��VPQ�M�Q�ҋu��P���%����M��=�����^��]� ����U����PL�EPQ���   �у�]� �U����PL�EP�EPQ�J�у�]� ���PL�BQ�Ѓ���������������̡��PL�BQ�Ѓ���������������̡��PL�BQ�Ѓ����������������U����PL�EP�EP�EPQ�J �у�]� ������������U����PL�EPQ��4  �у�]� �U����PL�EP�EP�EPQ�J$�у�]� ������������U����PL�EP�EP�EP�EPQ�J(�у�]� �������̡��PL�B,Q�Ѓ���������������̡��PL�B0Q�Ѓ����������������U����PL�EP�EPQ��  �у�]� ������������̡��PL���   Q�Ѓ�������������U����PL�E��  ��VPQ�M�Q�ҋu��P�������M�������^��]� ̡��PL�B4Q�Ѓ���������������̡��PL�B8j Q�Ѓ��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL�EPQ�J<�у�]� ���̡��PL�BQ��Y�U����PL�EP�EPQ�J@�у�]� U����PL�Ej PQ�JD�у�]� ��U����PL�Ej PQ�JH�у�]� ��U����PL�EjPQ�JD�у�]� ��U����PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��$���W�M�Q�U�R���������M����s����t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  �n���j�M�Q�U�R���}����M���r�������   ��U�R�Ѓ�^��]�����������U���$���UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}�����j�E�P�M�Q��������M��Qr�������   ��M�Q�҃�_^��]� ��U���$���UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��j��j�E�P�M�Q���y����M���q�������   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}����W�M�Q�U�R���������M����gq����t+�u�����������   ��U�R�Ѓ�_��^[��]� �����   �JL�E�P�ыu��P�����������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��D~��W�M�Q�U�R���4������M����p����t+�u������������   ��U�R�Ѓ�_��^[��]� �����   �JL�E�P�ыu��P���U��������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��}��W�M�Q�U�R���t������M�����o��_^��[t�����   ��U�R�������]Ë����   �J<�E�P���]������   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}���|��W�M�Q�U�R���ă�����M����7o����t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��$|��W�M�Q�U�R���������M����n����t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� �����̡��PL���   Q��Y��������������U����PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U����PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��z��W�M�Q�U�R��脁�����M�����l����t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���y��W�M�Q�U�R��贀�����M����'l����t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���x��W�M�Q�U�R���������M����Wk����t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��$x��W�M�Q�U�R��������M����j����t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  �ow��j�M�Q�UR���~~���M��i�������   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���v��j�U�R�E�P���~���M��fi�������   �
�E�P�у�^��]� ��������U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��zv��j�E�P�M�Q���}���M���h�������   ��M�Q�҃�_^��]� ��U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���u��j�E�P�M�Q���	}���M��ah�������   ��M�Q�҃�_^��]� ��U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��zu��j�E�P�M�Q���|���M���g�������   ��M�Q�҃�_^��]� ��U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���t��j�E�P�M�Q���	|���M��ag�������   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��t��j�U�R�E�P���{���M���f�������   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}��$t��W�M�Q�U�R���{�����M����f����t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��Ts��W�M�Q�U�R���Dz�����M����e����t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��r��W�M�Q�U�R���y�����M����e����t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��q��j�E�P�M�Q����x���M��!d�������   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��Oq��j�U�R�E�P���^x���M��c�������   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���p��j�U�R�E�P����w���M��Fc�������   �
�E�P�у�^��]� ��������U����H���   ]��������������U����H���   ]�������������̡��H���   ����H���   ��U����H���   V�u�R�Ѓ��    ^]�����������U����H���   ]��������������U����HL�QV�ҋ���u^]á��H�U�ER�UP���  RV�Ѓ���u���Q@�BV�Ѓ�3���^]����������U����H�U�E���  R�U�� P�ERP�у�]������U����H���   ]��������������U����H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡��PL�BLQ�Ѓ���������������̡��PL�BPQ�Ѓ����������������U����PL�EP�EPQ�JT�у�]� U����PL�EPQ��  �у�]� �U����PL�EPQ���   �у�]� ̡��PL�BXQ�Ѓ����������������U����PL�EP�EP�EPQ�J\�у�]� ������������U���4��SV��HL�QW�ҋ�3ۉ}�;��x  �M��������E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ����   �BSSW���Ѕ���   ���QL�BW�Ћ���;���   ��    �����   �B(���ЍM�Qh�   ���u�����������   �M�;���   �����   ���   S��;�tm�����   �ȋB<V�Ћ����   ���   �E�P�у�;�t���B@�HV�у���;��\����}��M�������M��I�����_^[��]� �}����B@�HW�ы����   ���   �M�Q�҃��M��y����M�����_^3�[��]� �����̡��PL�B`Q�Ѓ���������������̡��PL�BdQ�Ѓ����������������U����PL�EPQ�Jh�у�]� ���̡��PL��D  Q�Ѓ������������̡��PL�BlQ�Ѓ����������������U����PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Ehp� hP� h0� h � R�Q�U R�UR�UR�U���A�$�5��vLRP���   Q�Ѓ�4^]�  ������̡��PL���   Q�Ѓ�������������U����PL�EP�EP�EPQ��   �у�]� ���������U����PL��H  ]�������������̡��PL��L  ��U����PL��P  ]��������������U����PL��T  ]��������������U����PL�EP�EP�EP�EP�EPQ���   �у�]� �U����PL�EP�EP�EPQ���   �у�]� ���������U����PL�EP�EP�EP�EPQ��   �у�]� �����U����HL���   ]��������������U����HL���   ]��������������U����HL���   ]�������������̡��HL��  ����HL��@  ��h$�Ph^� �  ���������������U��Vh$�j\h^� ���Y  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� ��V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\���QLjP���   ���ЋM��U�Rh=���M�}��Ӫ���������   ���   �U�R�Ѓ��M��u�������_^��]Ë����   ���   �E�P�у��M��u��޾��_�   ^��]����U��� ��V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\���QLjP���   ���ЋM��U�Rh<���M�}������������   ���   �U�R�Ѓ��M��u��<�����_^��]Ë����   ���   �E�P�у��M��u�����_�   ^��]���̡�V�񋈈   ���   V�҃��    ^���������������U���EV���V��������Au���H��0  hxej,�����^��^]� �����U���W������G���U���d������A�  ������A��   ��e������AuR������AuKV��諘  ��褘  �ȅ�u��^����__��]Ëƙ����ʅ�u�u��E�^������__��]���������Au������=�e��������Au6�����������U������G�����_��������Au�����U����_�
����������]�  �E����U���e��������A{���������__��]�������������__��]����U����eV�E��������At����e������Au�������a����e�$�
�  �����a���^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3�����e;���W���$��葛  ��E����e�$�|�  �V����������Au���H��0  hxej�����^����_u������������^]� ���U������EV�ы�������z!���؋H��0  hxej5�����U������$��  �]��F�$�ۚ  �}��$�К  ��E�$�Ú  �^�����&���^��]� ��������������̋�� �e����������e���������̅�t��j�����̡��P��  ����P��(  ��U����P��   ��V�E�P�ҋuP��誻���M�������^��]� ��������̡��P��$  ��U����H��  ]��������������U����H���  ]�������������̡��H��  ��U����H���  ]��������������U����H��x  ]��������������U����H��|  ]��������������U���EV����et	V�X  ����^]� ��������������U��V�u���t���QP��Ѓ��    ^]���������̡��H��@  hﾭ���Y����������U��E��t���QP��@  �Ѓ�]����������������U����H���  ]��������������U����H��  ]�������������̡��H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW舙  ������u_^]Ã} tWj V�<�  ��_������F���   ^]���U����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW��  ������u_^]�Wj V�ƙ  ��_������F���   ^]�������������U����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW茘  ������u_^]�Wj V�F�  ��_������F���   ^]�������������U����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW��  ������u_^]�Wj V�Ƙ  ��_������F���   ^]�������������U����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW茗  ������u_^]�Wj V�F�  ��_������F���   ^]�������������U��M��t-�=�� t�y���A�uP�x�  ��]á��P�Q�Ѓ�]��������U��M��t-�=�� t�y���A�uP�8�  ��]á��P�Q�Ѓ�]��������U����H�U�R�Ѓ�]���������U����H�U�R�Ѓ�]���������U����E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�H�  ������u_^]�Wj V��  ��_������F���   ^]���������U����E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   ����t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�Y�  ������u_^]�Wj V��  ��_������F���   ^]����������U��E��w�   ����t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�Ɣ  ������u_^]�Wj V耕  ��_������F���   ^]�������U����H�U�R�Ѓ�]���������U����H�U�R�Ѓ�]���������U����H�U�R�Ѓ�]���������U����H�U�R�Ѓ�]���������U����Hp�]����Hp�h   �҃�������������U��V�u���t���QpP�B�Ѓ��    ^]���������U����Pp�EP�EPQ�J�у�]� U����Pp�EP�EPQ�J�у�]� U����Pp�EP�EPQ�J�у�]� U����Pp�EPQ�J�у�]� ����U����P�E���   ��VWP�EP�E�P�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ������������U��E��u� ��MP�EPQ�SL����]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h�ej;h0�j���������t
W���^����3��F��u_^]� �~ t3�9_��^]� ���H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ���H<�Q��3Ʌ����^��������������̃y t�   ËA��uË��R<P��JP�у��������U����u���H�]� ���J<�URP�A�Ѓ�]� ���������������U�� ���u���H�]Ë��J<�URP�A�Ѓ�]�U�� ���$V��u���H�1����J<�URP�A�Ѓ������Q�J�E�SP�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���[t.���B�u�HV�ы��B�P�M�Q�҃���^��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�u�QV�ҡ��H�A�U�VR�Ћ��Q�J�E�P�у���^��]���������������U�� ���$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�u�QV�ҡ��H�A�U�VR�Ћ��Q�J�E�P�у���^[��]����������������U�� ���$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у�����������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҋu�E�P��������Q�J�E�P�у���^[��]�������U�� ���$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h4fP�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у�����������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M���j h4f�M��B�����P�R@j �E�P�M�Q�M��҅����H�A�U�R���Ѓ���t/���Q�u�BV�Ћ��Q�J�E�P�у���^[��]Ë��M��B�PHjQ�M��ҡ��P�E�M��RLj�j�PQ�M��ҋu�E�P���k�����Q�J�E�P�у���^[��]���������������U����H<�A]����������������̡��H<�Q�����V��~ u>���t���Q<P�B�Ѓ��    W�~��t���ʧ��W�$������F    _^��������U���V�E�P���^�����P��������M��艧����^��]��̃=� uK� ���t���Q<P�B�Ѓ�� �    ����tV���@���V��������    ^������������U���8���H�AS�U�V3�R�]��Ћ��Q�JSj��E�h8fP�ы��B<�P�M�Q�ҋ���H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��T  �M�Q�U�R�M��hT  ����   W�}�}���   �����   �U��ATR�Ћ�����tB���Q�J�E�P���у��U�Rj�E�P���������Q�ȋBxW���E���t�E� ��t���Q�J�E�P����у���t���B�P�M�Q����҃��}� u"�E�P�M�Q�M��S  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3ۉ]�;�u_���H�A�U�R�Ћ��Q�JSj��E�h8fP�ы��B<�P�M�Q�ҋ���H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��R  �M�Q�U�R�M���R  ���p  W�}��I �E����   �����   �U��ATR�Ћ�������   ���Q�J�E�P���ы��B���   ���M�Qj�U�R���Ћ��Q�J���E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Bx��W�M����E��t�E ��t���Q�J�E�P����у���t���B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�����   P�BH�Ћ��Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��Q  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M���P  �EP�M�Q�M�u��u�-Q  ����   �u���E���tA��t<��uZ�����   �M�PHQ�ҋ��Q���ȋBxV�Ѕ�u-�   ^��]Ë����   �E�JTP��VP�[�������uӍUR�E�P�M��P  ��u�3�^��]����������V��~ u>���t���Q<P�B�Ѓ��    W�~��t��芢��W��������F    _^��������U��E�M�UP��P�EjP������]��������������̸   �����������U��V�u��t���u6�EjP��������u3�^]Ë�������t���t��U3�;P��I#�^]������̡��H\�������U����H\�AV�u�R�Ѓ��    ^]�������������̡��P\�BQ�Ѓ���������������̡��P\�BQ�Ѓ����������������U����P\�EPQ�J�у�]� ����U����P\�EP�EPQ�J�у�]� U����P\�EPQ�J�у�]� ���̡��P\�BQ�Ѓ����������������U����P\�EPQ�J �у�]� ����U����P\�EP�EPQ�J$�у�]� U����P\�EP�EP�EPQ�J(�у�]� ������������U����P\�EPQ�J0�у�]� ����U����P\�EPQ�J@�у�]� ����U����P\�EPQ�JD�у�]� ����U����P\�EPQ�JH�у�]� ���̡��P\�B4Q�Ѓ����������������U����P\�EP�EPQ�J8�у�]� U����P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu��F������H\�QV�҃���S���+���3���~=��I ���H\�U�R�U��EP�A(VR�ЋM��Q��������U�R������F;�|�_^[��]� ���������������U���VW�}�E��P���8����}� ��   ���Q\�BV�Ѓ��M�Q�������E���t]S3ۅ�~H�I �UR��������E�P�������E;E�!�����Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U��V�u�F��F�����������������|z  ����������D�Ez��^�P�P�]��������������N�X�N^�X]�������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��5�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A��e����������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E����X�X]� ��̋�3ɉ�H�H�H�V��V������FP�����3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  S�]���s  ��؋�U��M�U�>�U��@�����@�U��@�B�@�������@���@�   ;����U��p  �w�����  �w�������F�B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]؋�R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ʍU��R���[�[������E��KH��P�E�SL��H�щKP�P�ST�H�KX�P�����S\��z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����M��}������3�3����u��u�|+�A�����B�4�u�0u��u�p�����u�u�U�E;�}�Q���E����U��U��1���@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���@�D��KX�@�U�����]��C���@�K0���@�KH���C ��C�@�K8���@�KP���C(��C�C@�H���@3����KX���U��r  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������]��E�E����]���E����]��E׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���@�   �KXE)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� ����������h�Ph_� � ������������������h�jh_� ���������uË@����U��V�u�> t/h�jh_� ���������t��U�M�@R�Ѓ��    ^]���U��Vh�jh_� ����������t�@��t�MQ����^]� 3�^]� �������U��Vh�jh_� ���Y�������t�@��t�MQ����^]� 3�^]� �������U��Vh�jh_� ����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh�j h_� ����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh�j$h_� ���I�������t�@$��t�MQ����^]� 2�^]� �������Vh�j(h_� ����������t�@(��t��^��3�^������Vh�j,h_� �����������t�@,��t��^��3�^������U��Vh�j0h_� ����������t�@0��t�MQ����^]� 3�^]� �������U��Vh�j4h_� ���i�������t�@4��t�M�UQR����^]� ���^]� ��Vh�j8h_� ���,�������t�@8��t��^��3�^������U��Vh�j<h_� �����������t�@<��t�MQ����^]� ��������������U��Vh�j@h_� ����������t�@@��t�MQ����^]� ��������������U��Vh�jDh_� ���y�������t�@D��t�MQ����^]� 3�^]� �������U��Vh�jHh_� ���9�������t�@H��t�MQ����^]� ��������������Vh�jLh_� �����������t�@L��t��^��3�^������Vh�jPh_� �����������t�@P��t��^��3�^������Vh�jTh_� ����������t�@T��t��^��^��������Vh�jXh_� ���l�������t�@X��t��^��^��������Vh�j\h_� ���<�������t�@\��t��^��^��������U��Vh�j`h_� ���	�������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�jdh_� �����������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh�jhh_� ����������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh�jlh_� ���9�������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�jph_� �����������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh�jth_� ����������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�jxh_� ���i�������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh�j|h_� ���)�������t�@|��t�MQ����^]� 3�^]� �������U��Vh�h�   h_� �����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�h�   h_� ����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�h�   h_� ���6�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�h�   h_� �����������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������m�������_�U�^��[�U����U��������������������Xc  ����������D�Ez���P�P���]� �������E�����E����X�M��X��]� �������U���@�Pf�A���E�    �����]����]��]��Hf�������]����]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�����F�@��R�M��{����~���Q�M��i����v;�t�v��P�M��S����M����m��M�u�_^[�M�UQR�M�������]� ����������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$�h&�E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��&&+&?&S&����U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�����FP�~���3����F�F^��U��SV��WV�b����^S�Y����E3����~�~;�t_���Q���   hXf��jIP�у��;�t9�}��t;���B���   hXf��    jNQ�҃����uV�������_^3�[]� �E�~_�F^�   []� ����������U��SV��WV�����^S�����}3Ƀ��N�N;���   9��   �G;���   ���Q���  hXf��jlP�у����t=� t@�G��t9���JhXf��    ���  jqR�Ѓ����u���-���_^3�[]� �O�N�G�Q��    R�F�QP�]�������t�N�WP��QPR�h]����_^�   []� ���������U��SV��WV貿���~W詿��3Ƀ��N�N9M��   �E;���   ��    ���H���  hXfh�   S�҃����t=�} tH�E��tA���Q���  hXf��h�   P�у����u���2���_^3�[]� �U�V�,�F   ���H���  hXfh�   j�҃����t��E�M�F�PSPQ�a\���E����t!�V�?�W�RWP�E\����_^�   []� ��M�_^�   []� ���U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��S�]V��3�W�~���F�F�CV;C��   �����W����3��F�F���Q���   hXfjIj�Ѓ������   ���Q���   hXfjNj�Ѓ����uV薽����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� �P���W�J���3��F�F���B���   hXfjIj�у����t[���B���   hXfjNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP��������^]� ����������U��E��u�E�M�����   ]� �����������U��EHV����   �$�x-�   ^]á �@� ���uT�EP�W����=�.  }�����^]Ëu��t�h�fjmh0�j�˿������t ���u������tV���y���   ^]���    �   ^]ËM�UQR����������H^]�^]����- �u.�b����������t���,v��V膾������    �   ^]Ã��^]ÍI �,)-0-�,o--h$�Ph^� �������������������U��Vh$�jh^� ����������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �Vh$�jh^� ���L�������t�@��tV�Ѓ�^�3�^���U��Vh$�jh^� ����������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  Vh$�jh^� �����������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u���S����N`�K������   �@�����   �5�����ݞ�  ��^��]� ����U��Vh$�jh^� ���I�������t�@��t�M�UQRV�Ѓ�^]� ��������U��Vh$�jh^� ���	�������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��Vh$�j h^� �����������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh$�j$h^� ���y�������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��Vh$�j(h^� ���9�������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVh$�j,h^� �����������t �@,�E���t�E�MPQV�U���^��]� ��^��]� ��������U��Vh$�j0h^� ����������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������Vh$�j4h^� ���\�������t�@4��tV�Ѓ�^�3�^���Vh$�j8h^� ���,�������t�@8��tV�Ѓ�^�������U���`Vh$�jDh^� �����������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u���}�����^��]� ����U��Vh$�jHh^� ����������t�@H��t
�MQV�Ѓ�^]� ������������U��Vh$�jLh^� ���Y�������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��Vh$�jPh^� ����������t�@P��t
�MQV�Ѓ�^]� ������������U��Vh$�jTh^� �����������t�@T��t
�MQV�Ѓ�^]� ������������U��Vh$�jXh^� ����������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������Vh$�j`h^� ���<�������t�@`��tV�Ѓ�^�3�^���U��Vh$�jdh^� ���	�������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���Vh$�jhh^� �����������t1�@h��t*�MQ�U�VR�Ћu��P������M��	����^��]� �u���D	����^��]� �����������Vh$�jph^� ���\�������t�@p��tV�Ѓ�^Ã��^��Vh$�jlh^� ���,�������t�@l��tV�Ѓ�^Ã��^��Vh$�jth^� �����������t�@t��tV�Ѓ�^�3�^���U��Vh$�jxh^� �����������t�@x��t
�MQV�Ѓ�^]� ������������Vh$�j|h^� ����������t�@|��tV�Ѓ�^�������Vh$�h�   h^� ���Y�������t���   ��tV�Ѓ�^�U��Vh$�h�   h^� ���&�������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��Vh$�h�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���Vh$�h�   h^� ����������tU���   ��tKW�M�VQ�Ћ��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]� ���H�u�QV�҃���^��]� ����������Vh$�h�   h^� �����������t���   ��tV�Ѓ�^Ã��^������������U��Vh$�h�   h^� ����������t���   ��t
�MQV�Ѓ�^]� ������U��Vh$�h�   h^� ���f�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh$�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������Vh$�h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U��Vh$�h�   h^� ����������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��Vh$�h�   h^� ���6�������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��Vh$�h�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh$�h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh$�h�   h^� ���F�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh$�h�   h^� �����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������Vh$�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh$�h�   h^� ���i�������t���   ��tV�Ѓ�^�3�^�������������Vh$�h�   h^� ���)�������t���   ��tV�Ѓ�^�3�^�������������Vh$�h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U��Vh$�h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������Vh$�h�   h^� ���Y�������t���   ��tV�Ѓ�^�3�^�������������U���Vh$�h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh$�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh$�h�   h^� ���Y�������t���   ��tV�Ѓ�^�3�^�������������U���Vh$�h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh$�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh$�h�   h^� ���Y�������t���   ��tV�Ѓ�^�3�^�������������U��Vh$�h�   h^� ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVh$�h�   h^� �����������t#���   �E���t�E�MPQV�U���^��]� ��^��]� ��U��Vh$�h�   h^� ���v�������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��Vh$�h�   h^� ���&�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh$�h�   h^� �����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh$�h   h^� ����������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������Vh$�h  h^� ���9�������t��  ��tV�Ѓ�^�3�^�������������U���Vh$�h  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh$�h  h^� ���s�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh$�h  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��Vh$�h  h^� ���v�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh$�h  h^� ���6�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh$�h  h^� �����������t��  ��t
�MQV�Ѓ�^]� ������Vh$�h   h^� ��蹿������t��   ��tV�Ѓ�^�3�^�������������U��Vh$�h$  h^� ���v�������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh$�h(  h^� ���&�������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh$�h,  h^� ���־������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh$�h0  h^� ��艾������t��0  ��tV�Ѓ�^�3�^�������������U��Vh$�h4  h^� ���F�������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh$�h8  h^� �����������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh$�h<  h^� ��覽������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��Vh$�h@  h^� ���V�������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh$�hD  h^� ���	�������t��D  ��tV�Ѓ�^�3�^�������������U��Vh$�hH  h^� ���Ƽ������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh$�hL  h^� ���v�������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh$�hP  h^� ���&�������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVh$�hT  h^� ���ջ������t'��T  �E���t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��Vh$�hX  h^� ���v�������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��Vh$�j<h^� ���)�������t�@<��t�M�UQRV�Ѓ�^]� ��������U��Vh$�j@h^� ����������t�@@��t�MQV�Ѓ�^]� 3�^]� �����h(�Ph�� 谺�����������������h(�jh�� 菺������uË@����U��V�u�> t/h(�jh�� �c�������t��U�M�@R�Ѓ��    ^]���U��Vh(�jh�� ���)�������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh(�jh�� ���ٹ������t�@��t�M�UQR����^]� ����������U��Vh(�jh�� ��虹������t�@��t�M�UQR����^]� ����������U��Vh(�jh�� ���Y�������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh(�j h�� ���	�������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh(�j$h�� ��蹸������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh(�j(h�� ���i�������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh(�j,h�� ����������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��Vh(�j0h�� ��蹷������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh(�j4h�� ���i�������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVh(�j8h�� ����������t�@8�E���t�E�MPQ���U�^��]� ��^��]� ����������U��Vh(�j<h�� ��蹶������t�@<��t�M�UQR����^]� ����������U��Vh(�j@h�� ���y�������t�@@��t�M�UQR����^]� 3�^]� ���U��Vh(�jHh�� ���9�������t�@H��t�M�UQR����^]� 3�^]� ���U��Vh(�jDh�� �����������t�@D��t�M�UQR����^]� 3�^]� ���U��QVh(�jLh�� ��踵������t#�@L�E���t�E�EP�����$�U�^��]� ��^��]� �����U��Vh(�jPh�� ���i�������t�@P��t�M�UQR����^]� 3�^]� ���U��Vh(�jTh�� ���)�������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh(�jXh�� ���ٴ������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh(�j\h�� ��艴������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu h(�jh�� �2�������t�@�ЉF�~��t6h(�jh�� ��������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+h(�jh�� 豳������t�@��t�M�UQR���Ѓ~ t1h(�jh�� 耳������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u h(�jh�� �3�������t�@�ЉF�v��t+h(�jh�� ��������t�@��t�M�UQR����^]� �������������U��V�q��t@h(�jh�� �Ĳ������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<h(�j h�� �d�������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu h(�jh�� ��������t�@�ЉF�}�]�M�UWSQR���  ��t�N��t�E�UWSPR����_^[]� _^3�[]� �U��V�q��t8h(�j(h�� 褱������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��I��t)�E$�E�UP�E���\$�E�$R�UPR����]�  3�]�  �������U��V�q��t<h(�j0h�� ��������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U������   �BXQ�Ѓ���u]� ���Q|�M�RQ�MQP�҃�]� ���U������   �BXQ�Ѓ���u]� ���Q|�M�R8Q�MQP�҃�]� ���U��EV��j ����Qj j P�B�ЉF����^]� ��̡�Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ���Q�MP�EP�Q�JP�у��F�   ^]� ����U����PH�EPQ���  �у�]� �U����P�B4VW�}j��h�  ���ЋMWQ���D  _^]� ��������������U��V���PXW�ҋ}P���������Et�_�   ^]� �M�UPWQR���1  _^]� �����������U��S�]VW��j ���l����8�  �}uI�~ uC���P���   j h�  ���Ѕ�u���QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ����  _^[]� ��������U��EP�A    ������]� �����̸   �A� ������A   � ������U���@S�]VW����`��u�G   �}  ����   �M3�V�z����8�  u4����P�w蔏�����P�M�B4��jh�  ��_^�C�[��]� �MV�5����8�  u�E�M��RPQ����_^�   [��]� �MV�����8�  t�MV������8��  ���P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P譓��3��؃��u�;�t���QH���  VS�Ѓ��E��M�;O�f  9w�]  ���B�M���   Vh�  �҅�u!���P�M���   Vh�  �Ѕ��  ���Q�M�B4Vh�  ��;�t
V���������E��G�����   ���   �Ћ]�E�;���   ;���   S�7����M���jQ�ˉu��uĉuȉủuЉu؉u���r���U�E��ˉu��u�u�U�E��]��E�   ������t!��t��t�u���E�   ��E�   ��E�   �
7���M�;�t�N�����BX�M�Q����P��7���M܃�;�t�L����M��$L���M��L���M������]�M�U�EQSRP����  _^[��]� �M�����_^�   [��]� �������������̸   � ��������� ������������̃��� ����������� �������������U����H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� ���Q0�F�M���   PQW�ҋF��^_]� U����H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U����H���  ]��������������U����H���  ]��������������U����P�EP�EP�EP�EPQ���   �у�]� �����U����E�P�EP�E���\$�E�$PQ���   �у�]� �������������U����P�EP�EP�EPQ���   �у�]� ��������̡��P���   Q�Ѓ�������������U����P�EP�EP�EPQ���   �у�]� ���������U����P�EP�EPQ���   �у�]� �������������U����H�U�ApR�Ѓ�]� �����U����P�EP�EPQ���  �у�]� �������������U����P�EP�EPQ���  �у�]� �������������U����P�EP�EPQ���  �у�]� �������������U����P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P��)  ��R���E�P���ҡ��P�B<�M��Ћ}��t0j �M�QW��������u���B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4���@� �E��]�E� ^�E�`^�E��^�E��]�E��]�E�@^ǅx����^ǅ|����]�E�^�E�p^�E��]�E� ^�E��^�E��]�E��]�E�0^�E�P^�E��]�EĠ^�(0�������B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۉ]���u���H�A�UR�Ѓ�^3�[��]Ë��Q�B<W�M3��Ѕ��'  �\  �E���tq�MQ�M��	G��Wh�f�M�軴��P�M���F���u�Wj��U�R�E�P��\���Q�_?�Y����P��x���R�J����P�E�P�J����P���  �E���t�E� �� t�M�����G����t��x��������F����t��\��������F����t�M̃����F����t���Q�J�E�P����у���t�M��F���}� t"�U(�E$�M�R�UP�EQ�MRPQ���������U�R�O  ����E$�M�UVP�Ej QRP������������Q�J�EP�у���_^[��]����������������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`<����������̋�`L����������̋�`����������̋�` ����������̋�`0����������̋�`P����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`H����������̋�`����������̋�`����������̋�`,����������̡��H���   ��U����H���   V�u�R�Ѓ��    ^]����������̡��P���   Q�Ѓ�������������U����P�EPQ���   �у�]� ̡��H�������U����H�AV�u�R�Ѓ��    ^]��������������U����H�AV�u�R�Ѓ��    ^]��������������U����P��Vh�  Q���   �E�P�ы����   �Q8P�ҋ�����   ��U�R�Ѓ���^��]��������������̡��P�BQ�Ѓ����������������U����P�EPQ�J\�у�]� ����U����P�EP�EP�EP�EP�EPQ���   �у�]� �U����P�EP�EP�EP�EPQ�JX�у�]� �������̡��P�B Q��Y�U����P�EP�EP�EP�EPQ���   �у�]� �����U����P�EP�EP�EPQ�J�у�]� ������������U����H��   ]��������������U����P�R$]�����������������U����P�EP�EP�EP�EPQ�J(�у�]� ��������U����P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U����P�EP�EP�EP�EPQ�J,�у�]� ��������U���V��H�QWV�ҋ����H�QV�ҋ��Q�M�R4Q�MQ�MQOWHPj j V�҃�(_^]� ���������������U����P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U����P�EP�EPQ�J@�у�]� U����P�EPQ�JD�у�]� ���̡��P�BLQ�Ѓ���������������̡��P�BLQ�Ѓ���������������̡��P�BPQ�Ѓ����������������U����P�EPQ�JT�у�]� ����U����P�EPQ�JT�у�]� ����U����P�EP�EPQ���   �у�]� �������������U����P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �����   j P�BV�Ћ����   �
�E�P�у� ��^��]� ������̡��P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡��H�������U����H�AV�u�R�Ѓ��    ^]��������������U����P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U����P�EPQ�J�у�]� ���̡��P�BQ��Y�U����P�EP�EPQ�J�у�]� U��VW���ԁ���M�U�x@�EPQR��辁���H ���_^]� �U��VW��褁���M�U�xD�EPQR��莁���H ���_^]� �V���x����xH u3�^�W���f����΍xH�\����H �_^�����U��V���E����xL u3�^]� W���0����M�U�xL�EPQR�������H ���_^]� �������������U��V��������xP u���^]� W���߀���M�U�xP�EP�EQRP���ŀ���H ���_^]� ��������U��V��襀���xT u���^]� W��菀���M�xT�EPQ���}����H ���_^]� U���S�]VW���t.�M���Y�����O����xL�E�P���A����H ��ҍM��0Z���}��tZ���H�A�U�R�Ћ��Q�J�E�WP�ы��B�P�M�Q�҃��������@@��t���QWP�B�Ѓ�_^[��]� ������U��VW������xH�EP������H ���_^]� ���������U��VW������M�U�xD�EP�EQRP���j���H ���_^]� �������������U��V���E���xP u
�����^]� W���-���M�U�xP�EP�EQ�MR�UPQR������H ���_^]� ��������������U��V����~���xT u
�����^]� W����~���M�xT�EPQ���~���H ���_^]� ��������������U��V���~���xX tW���~���xX�EP���y~���H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��  ����t.�E�;�t'���J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡��H��   ��U����H��$  V�u�R�Ѓ��    ^]�����������U����UV��H��(  VR�Ѓ���^]� �����������U����P�EQ��,  P�у�]� �U����P�EQ��,  P�у����@]� �����������̡��H��0  ����H��4  ��U��E��t�@�3����RP��8  Q�Ѓ�]� �����U����P�EPQ��<  �у�]� �U����P�EP�EP�EPQ��@  �у�]� ���������U����P�EP�EPQ��D  �у�]� �������������U����P�EPQ��H  �у�]� �U����P�E��L  ��VWPQ�M�Q�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ��������������̡��P��T  Q�Ѓ������������̡��P��P  Q�Ѓ�������������U����P�EPQ��X  �у�]� ̡��H��\  ��U����H��`  V�u�R�Ѓ��    ^]�����������U����P�EP�EP�EP�EP�EPQ��d  �у�]� �U����P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w���6����3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7���Oz���xP t$S���Az��j j �XPj�FP���-z���H ���[�    �~` t���H�V`�AR�Ѓ��F`    _^������������U��SV��Fx���Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR�d"������u#���h�f���H��0  h�   �҃��E�~P���8���j j jW�N����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ���Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ������F|��u�E�~x��t�    �F`_^]� �M�Fx������t�3�_^]� U��QVW�}����>  ���H�QhV�҃�����u"�H��0  h�fh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���  �EF;u�|�UR�y����_�   ^��]� �������������U��QVW�}����~  ���H�QhV�҃�����u"�H��0  h�fh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'�����QP�Bh�Ѓ���t�M��R���,  F;u�|ʍEP�-x����_�   ^��]� �������������h�fh�   h0�h�   ��{������t�������3��������V���(����N^�2�����������������U��VW�}�7��t��������N�2��V��z�����    _^]�h,�Ph�f �0������������������U��h,�jh�f ��������t
�@��t]�����]�������U��Vh,�jh�f �ۏ��������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�1���E�NP�у�4�M����1����^]ÍM�1�����^]��U��h,�jh�f �l�������t
�@��t]��3�]��������U��h,�jh�f �<�������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^á��H�F��  h8gj8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� }(�V;Vu��������t�F�N��    �F9~|؋V;Vu���������t��F�N�U���F_�   ^]� ��������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T����H;ǉ�F�M���F_�   ^]� ����U��E��|2�Q;�}+J;Q}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�St��3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W��g�]r��3����_�F�F^��������������U���SV�uW���^S�}��&r��3���F�F�O�N�W���V9G�E~|��I �O���F�U�9FuL��u�~��~��t���< ��tY���H���  h8gj8��    RP�у���t0�~�}���V��M����E�F@;G�E|�_^�   [��]� _^3�[��]� U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|���P�����_^]� �U����E�Qj�E��ARP�M��E��g�+�����]� �����U����Q�Ej�E��A�MRPQ�M��E��g�G�����]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q�0g��t!�A��t�B�A�Q�P�A    �A    �̋�� �g�@0g�HV3��q�q�P�r�r�0g�p�p�p�P�H^������V����g�����F3��F0g;�t�N;�t�H�F�N�H�V�V�F�F0g;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3��0g;�t�F;�t�A�F�N�H�V�V�Et	V�r������^]� ������������U��V��W�~W��g�n��3����E��F�Ft	V��q����_��^]� ������U��V��������Et	V�q������^]� �I��8��<�0��@���D���H����L��P����T����X���\���Ë�U�������F  �} �8�t��  ��]�;��u���L  ��U��EVW��u|P�*  Y��u3��  �  ��u�*  ���%*  �`�T���(  �@���"  ��}�#  ���	(  ��| �%  ��|j �   Y��u�<��   �%  ��3�;�u19=<�~��<�9=��u�F"  9}u{��$  ��  �*  �j��uY�|  h  j��  ��YY;��6���V�5`��5|���  Y�Ѕ�tWV�  YY�`�N���V�  Y�������uW�7  Y3�@_^]� jh���+  ����]3�@�E��u9<���   �e� ;�t��u.��g��tWVS�ЉE�}� ��   WVS�r����E����   WVS�̯���E��u$��u WPS踯��Wj S�B�����g��tWj S�Ѕ�t��u&WVS�"�����u!E�}� t��g��tWVS�ЉE��E������E���E��	PQ�*  YYËe��E�����3���*  Ë�U��}u�~,  �u�M�U�����Y]� ��������������̃=(� t-U�������$�,$�Ã=(� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�Ë�Q��g��,  YË�U��V��������EtV��m��Y��^]� ����U��WV�u�M�}�����;�v;���  ��   r�=(� tWV����;�^_u^_]�"1  ��   u������r*��$����Ǻ   ��r����$��~�$����$���~�~�~#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I {h`XPH@8�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$� ������$�Ѐ�I �Ǻ   ��r��+��$�$��$� ��4�X����F#шG��������r�����$� ��I �F#шG�F���G������r�����$� ���F#шG�F�G�F���G�������V�������$� ��I Ԁ܀��������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$� ���0�8�H�\��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̺��!0  ���/  �Ƀ=8�t�����=  �����z�����������������̃= � �D  ���\$�D$%�  =�  u�<$f�$f��f���d$��C  � �~D$f(�gf(�f(�fs�4f~�fT�gf��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�@  ���D$��~D$f��f(�f��=�  |!=2  �fT�g�\�f�L$�D$����f��gfV�gfT�gf�\$�D$�jhІ�$  �e� �u;5�w"j�E  Y�e� V�$M  Y�E��E������	   �E��$  �j�D  YË�U��V�u�����   SW�=`�=̻ u�R+  j�)  h�   �*  YY�0���u��t���3�@P���uV�S���Y��u��uF�����Vj �5̻�׋؅�u.j^9X�t�u��O  Y��t�u�{����O  �0�~O  �0_��[�V��O  Y�jO  �    3�^]������̋T$�L$��ti3��D$��u��   r�=(� t�P  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh���#  �u��tu�=0�uCj�C  Y�e� V�C  Y�E��t	VP��C  YY�E������   �}� u7�u�
j�oB  Y�Vj �5̻�`��u�hN  ���`P�N  �Y��"  Ë�U��QSVW�5H��  �5D����}��t  ��YY;���   ��+ߍC��rwW�uO  ���CY;�sH�   ;�s���;�rP�u��S  YY��u�G;�r@P�u��=  YY��t1��P�4��  Y�H��u�  ���V�v  Y�D��EY�3�_^[�Ë�Vjj �  ��V�O  ���H��D���ujX^Ã& 3�^�jh��!  �  �e� �u�����Y�E��E������	   �E��!  ��  Ë�U���u���������YH]����������̃��$��O  �   ��ÍT$�O  R��<$�D$tQf�<$t�`O  �   �u���=4� ��O  �   �0���O  �  �u,��� u%�|$ u���5O  �"��� u�|$ u�%   �t����-���   �=4� �vO  �   �0��N  ZË�U��EV���F ��uc��  �F�Hl��Hh�N�;ȭt���Hpu��Y  ��F;�t�F���Hpu�IR  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P��\  ��e�F�P�[  ��Yu��P�\  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P��[  �M��E��M��H��EP�\  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�s`  @PV�V��\  ��^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M�������3�;�u+��I  j_VVVVV�8�WY  ���}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�I  j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h hSV��_  ��3ۅ�tSSSSS�hW  ���N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F���t�90uj�APQ�u[  ���}� t�E��`p�3�_^[�Ë�U���,���3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�a  3ۃ�;�u�hH  SSSSS�0��W  �����o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q�$_  ��;�t���u�E�SP�u��V�u��������M�_^3�[�D����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �C���9}}�}�u;�u+�~G  j^WWWWW�0��V  ���}� t�E�`p����  9}vЋE��� 9Ew	�@G  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�J  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� ��_  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �y_  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�������u�E�8 u���} �4����$�p���WF�_  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP��]  0�F�U�����;�u��|��drj jdRP�]  0��U�F����;�u��|��
rj j
RP�]  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N�������u-�D  j^�03�PPPPP�S  ���}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V�������}� t�E��`p�3�_^[�Ë�U���,���3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�[  3ۃ�;�u�C  SSSSS�0�uR  �����Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P��Y  ��;�t���u�E�SV�u���`������M�_^3�[������Ë�U���0���3ŉE��ESV�uWj_W�M�Q�M�Q�p�0��Z  3ۃ�;�u�SB  SSSSS�8�Q  �����   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW�$Y  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[�����Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3���8��6�  ��Y���(r�_^Ë�Vh   h   3�V��Z  ����tVVVVV��N  ��^Ë�U����h�]��h�]��E��u��M��m��]����]�����z3�@��3���h4h�`��thhP�`��tj ���������U���(  �X��T��P��L��5H��=D�f�p�f�d�f�@�f�<�f�%8�f�-4���h��E �\��E�`��E�l����������  �`��\��P�	 ��T�   �������������������0`���j�Z  Yj �,`h@h�(`�=�� uj��Y  Yh	 ��$`P� `�Ë�U��V�5d��58`�օ�t!�`����tP�5d����Ѕ�t���  �'�XhV�4`��uV�  Y��thHhP�`��t�u�ЉE�E^]�j ����YË�U��V�5d��58`�օ�t!�`����tP�5d����Ѕ�t���  �'�XhV�4`��uV�   Y��ththP�`��t�u�ЉE�E^]��<`� ��V�5d��8`����u�5x��e���Y��V�5d��@`��^á`����tP�5���;���Y�Ѓ`���d����tP�D`�d���c1  jh0��  �XhV�4`��uV�a  Y�E�u�F\�h3�G�~��t$hHhP�`�Ӊ��  hth�u��Ӊ��  �~pƆ�   CƆK  C�Fh��j�2  Y�e� �vh�H`�E������>   j��1  Y�}��E�Fl��u�ȭ�Fl�vl�qI  Y�E������   �  �3�G�uj��0  Y�j��0  YË�VW�`�5`��������Ћ���uNh  j��  ��YY��t:V�5`��5|������Y�Ѕ�tj V�����YY�`�N���	V����Y3�W�L`_��^Ë�V��������uj�>  Y��^�jhX��  �u����   �F$��tP�P���Y�F,��tP�B���Y�F4��tP�4���Y�F<��tP�&���Y�F@��tP����Y�FD��tP�
���Y�FH��tP�����Y�F\=�htP�����Yj�0  Y�e� �~h��tW�P`��u����tW����Y�E������W   j�P0  Y�E�   �~l��t#W�cH  Y;=ȭt���t�? uW�oF  Y�E������   V�f���Y��  � �uj�/  YËuj�/  YË�U��=`��tK�} u'V�5d��58`�օ�t�5`��5d����ЉE^j �5`��5|�����Y���u�x����d����t	j P�@`]Ë�VW�XhV�4`��uV�R  Y�����^  �5`h�hW��h�hW�t���h�hW�x���h�hW�|��փ=t� �5@`���t�=x� t�=|� t��u$�8`�x��D`�t���5|�����<`�d������   �5x�P�օ���   �_  �5t������5x��t������5|��x������5���|��u����������,  ��teh��5t������Y�У`����tHh  j�   ��YY��t4V�5`��5|�����Y�Ѕ�tj V�y���YY�`�N��3�@��$���3�_^Ë�U��VW3��u�������Y��u'9��vV�T`���  ;��v��������uʋ�_^]Ë�U��VW3�j �u�u�qS  ������u'9��vV�T`���  ;��v��������uË�_^]Ë�U��VW3��u�u�ET  ��YY��u,9Et'9��vV�T`���  ;��v��������u���_^]Ë�U��W��  W�T`�u�4`���  ��`�  w��t�_]Ë�U���a  �u�  �5h��D���h�   �Ѓ�]Ë�U��h�h�4`��th�hP�`��t�u��]Ë�U���u�����Y�u�X`�j�n,  Y�j�+  YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=�g th�g�U  Y��t
�u��gY�B���hDah,a����YY��uBhT������� a�$(a�c����=P� YthP��bU  Y��tj jj �P�3�]�jh���  j�+  Y�e� 3�C9����   ����E����} ��   �5H������Y���}؅�tx�5D�����Y���u܉}�u����u�;�rW����9t�;�rJ�6��������������5H��~������5D��q�����9}�u9E�t�}�}؉E����u܋}��hTa�Ha�_���Yh\a�Xa�O���Y�E������   �} u(���j�)  Y�u�����3�C�} tj�)  Y��7
  Ë�U��j j�u�������]�jj j ������Ë�V������V�5  V�W  V�C  V��  V��V  V��T  V�  V�T  h��������$�h�^�jTh���r	  3��}��E�P�h`�E�����j@j ^V�&���YY;��  �@��54���   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@�@���   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M���@���4� ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=4�|���=4��e� ��~m�E����tV���tQ��tK�uQ�d`��t<�u���������4�@��E� ���Fh�  �FP�mU  YY����   �F�E�C�E�9}�|�3ۋ���5@�����t���t�N��r�F���uj�X�
��H������P�``�����tC��t?W�d`��t4�>%�   ��u�N@�	��u�Nh�  �FP��T  YY��t7�F�
�N@�����C���g����54��\`3��3�@Ëe��E���������p  Ë�VW�@��>��t1��   �� t
�GP�l`���@   ;�r��6������& Y����@�|�_^Ã=L� u�=  V�5@�W3���u����   <=tGV�H  Y�t���u�jGW�n�����YY�=����tˋ5@�S�BV�\H  ��C�>=Yt1jS�@���YY���tNVSP��H  ����t3�PPPPP�L@  �����> u��5@��
����%@� �' �@�   3�Y[_^��5��������%�� ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�S  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#��R  Y��t��M�E�F��M��E���R  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9L�u��:  h  ���VS�Ļ�p`�T��5��;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�q�����Y;�t)�U��E�P�WV�}�������E���H����5��3�����_^[�Ë�U��Ȼ��SV�5�`W3�3�;�u.�֋�;�t�Ȼ   �#�`��xu
jX�Ȼ��Ȼ����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5�`SSS+�S��@PWSS�E��։E�;�t/P����Y�E�;�t!SS�u�P�u�WSS�օ�u�u�����Y�]��]�W�|`���\��t;�u��x`��;��r���8t
@8u�@8u�+�@P�E��0�����Y;�uV�t`�E����u�VW�������V�t`��_^[�Ë�V������W��;�s���t�Ѓ�;�r�_^Ë�V������W��;�s���t�Ѓ�;�r�_^Ë�U��3�9Ej ��h   P��`�̻��u]�3�@�0�]Ã=0�uWS3�9�W�=`~3V�5���h �  j �v���`�6j �5̻�׃�C;�|�^�5�j �5̻��_[�5̻��`�%̻ �Ë�U��QQV�G��������F  �V\���W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ����=�����;�}$k��~\�d9 �=�����B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]��h �d�5    �D$�l$�l$+�SVW���1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35��W��E� �E�   �{���t�N�38�����N�F�38�{����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���8N  �E���|@G�E��؃��u΀}� t$����t�N�38�����N�V�3:������E�_^[��]��E�    �ɋM�9csm�u)�=,� t h,���H  ����t�UjR�,����M��M  �E9Xth��W�Ӌ���M  �E�M��H����t�N�38�u����N�V�3:�e����E��H���qM  �����9S�R���h��W���M  ������U�������e� �e� SW�N�@��  ��;�t��t	�У���`V�E�P��`�u�3u���`3��`3���`3��E�P��`�E�3E�3�;�u�O�@����u������5���։5��^_[��jh���r����e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E��t���Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[�������(�3��jh������j�,  Y�e� �u�N��t/�Ի�л�E��t9u,�H�JP�V���Y�v�M���Y�f �E������
   ����Ë���j��  Y���������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�U���(  ���3ŉE��ТVtj
��   Y�G  ��tj�G  Y�Т��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P�I�������������(�����0���j ǅ����  @��������,����,`��(���P�(`j����̋�U��QQS�]VW3�3��}�;�آt	G�}���r���w  j�L  Y���4  j�sL  Y��u�=L��  ���   �A  h�n�  S�ػW�<  ����tVVVVV�4  ��h  ��Vj ��� �p`��u&h�nh�  V�O<  ����t3�PPPPP��3  ��V�;  @Y��<v8V�;  ��;�j��h�n+�QP�K  ����t3�VVVVV�3  ���3�h�nSW�kJ  ����tVVVVV�n3  ���E��4�ܢSW�FJ  ����tVVVVV�I3  ��h  h�nW�H  ���2j��``��;�t$���tj �E�P�4�ܢ�6��:  YP�6S��`_^[��j�K  Y��tj��J  Y��u�=L�uh�   �)���h�   ����YYË�U��E���]�U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ë�U��� S3�9]u ��"  SSSSS�    �K2  ������   �MV�u;�t!;�u�"  SSSSS�    �2  ������S�����E�;�w�M�W�u�E��u�E�B   �u�u�P�u��GK  ����;�t�M�x�E����E�PS�I  YY��_^[�Ë�U���uj �u�u�u�5�����]�����U���0���S�ٽ\�����=� t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=� t�#  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����,  �   [�À�8�����=4� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �8o�����������(o����s4�Ho�,ǅr���   �0o����������� o����v�@oVW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�T  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����D   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Àzuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp���������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-����p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t��������� u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t�У���У���l$����ԣ���ԣ���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r �������أ�|$�l$�ɛ�l$������l$��Ã�,��?�$������,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  ������ܣ �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�������Ƀ�u�\$0�|$(���l$�-������l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8����l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w������|$����<$� �|$$�D$$   �D$(�l$(������<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  ������ܣ �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�������Ƀ�u�\$0�|$(���l$�-������l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8����l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w������|$����<$� �|$$�D$$   �D$(�l$(������<$�l$$�Q�����0Z�����0Z�������@���������Ë�U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9��t�5$��T���Y��	�M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E�p��M��]�Q��]���]���Y����  �z  � "   �  �E�p��M��]�Q��E�   �]���]���Y�j  �E�   �E�p��E� p��]���]���"  �M��E� p�r����E��o�׉M��E��o�Z����E�p놃�tNIt?It0It ��t����   �E��o��E��o��E�p����E�p�x����E�   ��������   �E�   �E��o��������������   �$����E��o��E� p��E�p��E��o��E��o��E��o�y����E��o�m����E��o��Eܼo��Eܸo��M����]���]�M��]�Q�E�   ��Y��u��  � !   �E��_^[������ �	�����'�����3�<�E��% � ����� �3�Ë�U��QQSV���  V�5 ��K  �EYY�M�ظ�  #�QQ�$f;�uU�?J  YY��~-��~��u#�ESQQ�$j��H  ���rVS�MK  �EYY�d�ES��a���\$�E�$jj�?�I  �]��EY�]�Y����DzVS�K  �E�YY�"�� u��E�S���\$�E�$jj�H  ��^[�Ë�VW3�� ��<�,�u��(��8h�  �0���6.  YY��tF��$|�3�@_^Ã$�(� 3����S�l`V�(�W�>��t�~tW��W�f����& Y����H�|ܾ(�_���t	�~uP�Ӄ���H�|�^[Ë�U��E�4�(���`]�jh ��7���3�G�}�3�9̻u�,���j�z���h�   ����YY�u�4�(�9t���nj����Y��;�u�  �    3��Qj
�Y   Y�]�9u,h�  W�--  YY��uW蔼��Y�m  �    �]���>�W�y���Y�E������	   �E�������j
�(���YË�U��EV�4�(��> uP�"���Y��uj�����Y�6��`^]Ë�U�����k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �P�����   ���5�`h @  ��H� �  SQ�֋��P��   ���	P�P��@������    �P��@�HC�P��H�yC u	�`��P��x�ueSj �p�֡P��pj �5̻�`���P�k���+ȍL�Q�HQP�  �E����;P�v�m�����E�P��=�[_^�á�V�5�W3�;�u4��k�P�5�W�5̻��`;�u3��x���5���k�5�h�A  j�5̻�`�F;�t�jh    h   W��`�F;�u�vW�5̻�`뛃N��>�~���F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W��`��u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U������Mk��������M���SI�� VW}�����M���������3���U�������S�;#U�#��u
���];�r�;�u����S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1���	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t���C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;P�u�M�;�u�%P� �M���B_^[�Ë�U��E3�;�H�tA��-r�H��wjX]Ë�L�]�D���jY;��#���]�������u���Ã��������u���Ã�Ë�U��V������MQ�����Y�������0^]Ë�U��E�T�]Ë�U���5T������Y��t�u��Y��t3�@]�3�]�U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh ������3��]3�;���;�u�y����    WWWWW��  ������S�=0�u8j����Y�}�S�A���Y�E�;�t�s���	�u���u��E������%   9}�uSW�5̻��`���������3��]�u�j�����Y���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�2  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��p�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��<p�����������,p�����   s��Lp��4p�����������$p�����   v��Dp�����U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�-���3��ȋ��~�~�~����~���������F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  ���3ŉE�SW������P�v��`�   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R�j�����C�C��u�j �v�������vPW������Pjj �X?  3�S�v������WPW������PW�vS�9=  ��DS�v������WPW������Ph   �vS�=  ��$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[������jh@�������(��������Gpt�l t�wh��uj �[���Y��������j�,���Y�e� �wh�u�;5�t6��tV�P`��u����tV�V���Y���Gh�5��u�V�H`�E������   뎋u�j�����YË�U���S3�S�M�蟬���\����u�\�   ��`8]�tE�M��ap��<���u�\�   ��`�ۃ��u�E��@�\�   ��8]�t�E��`p���[�Ë�U��� ���3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9����   �E��0=�   r����  �p  ����  �d  ��P��`���R  �E�PW��`���3  h  �CVP芨��3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�C����M��k�0�u��� ��u��*�F��t(�>����E����D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C����Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95\��X�������M�_^3�[������jh`�������M���������}�������_h�u�u����E;C�W  h   �8���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�P`��u�Fh=��tP�2���Y�^hS�=H`���Fp��   ����   j����Y�e� �C�l��C�p��C�t�3��E��}f�LCf�E`�@��3��E�=  }�L���@��3��E�=   }��  ���@���5��P`��u��=��tP�y���Y��S���E������   �0j�&���Y��%���u ����tS�C���Y�����    ��e� �E�����Ã=L� uj��V���Y�L�   3�Ë�U��SV�u���   3�W;�to=�th���   ;�t^9uZ���   ;�t9uP�ʥ�����   �z;  YY���   ;�t9uP詥�����   �;  YY���   葥�����   膥��YY���   ;�tD9u@���   -�   P�e������   ��   +�P�R������   +�P�D������   �9��������   �=(�t9��   uP��8  �7����YY�~P�E   ���t�;�t9uP����Y9_�t�G;�t9uP�֤��Y���Mu�V�Ǥ��Y_^[]Ë�U��SV�5H`W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5P`W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Å�t7��t3V�0;�t(W�8�����Y��tV�E����> Yu���tV�Y���Y��^�3��jh���u���輵������Fpt"�~l t襵���pl��uj ����Y�������j����Y�e� �Fl�=ȭ�i����E��E������   ��j����Y�u�Ë�U��E���]Ë�U���(  ���3ŉE������� SjL������j P�/�����������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������0`j ���,`��(���P�(`��u��uj�H  Yh ��$`P� `�M�3�[������Ë�U���5���ı��Y��t]��j�	  Y]������U����u�M������E����   ~�E�Pj�u�A8  ������   �M�H���}� t�M��ap��Ë�U��=x� u�E����A��]�j �u����YY]Ë�U���SV�u�M�脣���]�   ;�sT�M胹�   ~�E�PjS�7  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�8  YY��t�Ej�E��]��E� Y��1���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P��1  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=x� u�E�H���w�� ]�j �u�����YY]Ë�U���(���3ŉE�SV�uW�u�}�M��2����E�P3�SSSSW�E�P�E�P��A  �E�E�VP�f7  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�l����Ë�U���(���3ŉE�SV�uW�u�}�M�芡���E�P3�SSSSW�E�P�E�P�SA  �E�E�VP�<  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�Ĕ������������������U��WV�u�M�}�����;�v;���  ��   r�=(� tWV����;�^_u^_]�"�����   u������r*��$�����Ǻ   ��r����$����$�����$���������#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I {�h�`�X�P�H�@�8��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$� ������$����I �Ǻ   ��r��+��$�$��$� ��4�X����F#шG��������r�����$� ��I �F#шG�F���G������r�����$� ���F#шG�F�G�F���G�������V�������$� ��I ���������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$� ���0�8�H�\��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��MS3�VW;�t�};�w�1���j^�0SSSSS���������0�u;�u��ڋъ�BF:�tOu�;�u������j"Y�����3�_^[]Ë�U��MSV�u3�W�y;�u�����j^�0SSSSS�.��������   9]v݋U;ӈ~���3�@9Ew����j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�a���@PWV�������3�_^[]Ë�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���H���u��P������Ɂ���  �P���t�M�_^f�H[�Ë�U���0���3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��A  �uЉC�E։�EԉC�E�P�uV������$��t3�PPPPP�<������M�_�s^��3�[�G������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j蹭��YË�U��E�M%����#�V������t1W�}3�;�tVV�J  YY�����j_VVVVV�8� �������_��uP�u��t	�QJ  ���HJ  YY3�^]Ã%� �jh��蘹���M3�;�v.j�X3���;E�@u�4����    WWWWW������3���   �M��u;�u3�F3ۉ]���wi�=0�uK������u�E;�w7j����Y�}��u����Y�E��E������_   �]�;�t�uWS�V�����;�uaVj�5̻�`��;�uL9=X�t3V�����Y���r����E;��P����    �E���3��uj�G���Y�;�u�E;�t�    ���̸���jh���z����]��u�u�����Y��  �u��uS�2���Y�  �=0���  3��}�����  j����Y�}�S�����Y�E�;���   ;5�wIVSP��������t�]��5V����Y�E�;�t'�C�H;�r��PS�u��L���S�����E�SP������9}�uH;�u3�F�u������uVW�5̻�`�E�;�t �C�H;�r��PS�u������S�u��b������E������.   �}� u1��uF������uVSj �5̻��`����u�]j�����YË}����   9=X�t,V�1���Y������������9}�ul���`P�v���Y��_����   ����9}�th�    �q��uFVSj �5̻��`����uV9X�t4V�����Y��t���v�V����Y�Z����    3��ٶ����G����|�����u�9������`P������Y��������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h��h �d�    P��SVW���1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh ������N����@x��t�e� ���3�@Ëe��E������(���� ����h���U���Y���Ë�U��E������������]Ë�U��E���V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5���i���Y�j h ��[���3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�������}؅�u����a  �������`�w\���]���������Z�Ã�t<��t+Ht�����    3�PPPPP������뮾�������������
�������E�   P襠���E�Y3��}���   9E�uj蘩��9E�tP�����Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.����M܋������9M�}�M�k��W\�D�E���������E������   ��u�wdS�U�Y��]�}؃}� tj ����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3������Ë�U��E���]Ë�U��E���]�jh@�荲���e� �u�u��`�E��/�E� � �E�3�=  �����Ëe�}�  �uj�L`�e� �E������E�����Ë�U����u�M�萑���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]���SVW�T$�D$�L$URPQQhd�d�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�F  �   �C�$F  �d�    ��_^[ËL$�A   �   t3�D$�H3��@���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�oE  3�3�3�3�3���U��SVWj j h�Q�e  _^[]�U�l$RQ�t$������]� ��U���SVW�`����e� �= � ����   h\x��`�����*  �5`hPxW�օ��  P誜���$@xW� ���P蕜���$,xW����P耜���$xW����P�k���Y����th�wW��P�S���Y����;�tO9�tGP豜���5���褜��YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9��;�t0P�a���Y��t%�ЉE���t��;�tP�D���Y��t�u��ЉE��5 ��,���Y��t�u�u�u�u����3�_^[�Ë�U��ES3�VW;�t�};�w����j^�0SSSSS���������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��e���j"Y����3�_^[]Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w�#���j^�0SSSSS����������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x��������j"Y���낋�U��MV3�;�|��~��u�H��(�H��H���n���VVVVV�    ����������^]Ë�U��E��t���8��  uP�Y���Y]Ë�U��QV�uV�wO  �E�FY��u����� 	   �N ����/  �@t������ "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�TM  �� ;�t�HM  ��@;�u�u��L  Y��uV�L  Y�F  W��   �F�>�H��N+�I;��N~WP�u�uK  ���E��M�� �F����y�M���t���t�����������@���p��@ tjSSQ��B  #����t%�F�M��3�GW�EP�u�K  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u�C����8*u�ϰ?�d����} �^[]Ë�U���x  ���3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������u�����u5�����    3�PPPPP������������ t
�������`p������
  �F@u^V��L  Y�p����t���t�ȃ��������@�����A$u����t���t�ȃ������@�����@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw����`x��3��3�3�����xj��Y������;���	  �$����������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�������Q  Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u��������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P��I  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ��������P����Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7���������{G  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V�+���������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5P��$���Y�Ћ���������   t 9�����u������PS�5\������Y��YY������gu;�u������PS�5X��А��Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�I7  ��0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u���������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF�D  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t�������*}�������� Y���������������t������������������������� t
�������`p��������M�_^3�[�!s���Ð������@������� ��S��QQ�����U�k�l$���   ���3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�(  ��h��  ��x����  �>YYt�=� uV�    Y��u�6��  Y�M�_3�^��q����]��[�3�Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u��`�M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M�������{L�H��M�����{,���2��M�����z�����M�����z�خ��خ��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E����a�S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�X���� "   ]��K���� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3����;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�U�������uV�,���Y�E�^�Ë����h��  �u(�  �u�����E ���Ë�U��=� u(�u�E���\$���\$�E�$�uj�/�����$]��4���h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   ���3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=� u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3���j����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�- ��]���t����- ��]�������t
�-��]����t	�������؛�� t���]����jh`�葕��3�9(�tV�E@tH9�t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%� �e��U�E�������e��U�q���Ë�U������3ŉE�SV3�W��9�u8SS3�GWhTyh   S��`��t�=���`��xu
��   9]~"�M�EI8t@;�u�����E+�H;E}@�E������  ;���  ����  �]�9] u��@�E �5�`3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�*  ��;�t� ��  �P�o��Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5�`SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�B)  ��;�tj���  ���P��n��Y;�t	� ��  �����3�;�tA�u�VW�u��u�u��`��t"SS9]uSS��u�u�u�VS�u ��`�E�V�g���Y�u��^����E�Y�Y  �]�]�9]u��@�E9] u��@�E �u�6  Y�E���u3��!  ;E ��   SS�MQ�uP�u ��6  ���E�;�tԋ5�`SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�,(  ��;�t����  ���P��m��Y;�t	� ��  �����3�;�t��u�SW�n�����u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��6  ���u������#u�W�<���Y��u�u�u�u�u�u��`��9]�t	�u��n��Y�E�;�t9EtP�un��Y�ƍe�_^[�M�3��d���Ë�U����u�M���p���u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap��Ë�U��QQ���3ŉE���SV3�W��;�u:�E�P3�FVhTyV��`��t�5��4�`��xu
jX���������   ;���   ����   �]�9]u��@�E�5�`3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�E&  ��;�t� ��  �P��k��Y;�t	� ��  ���؅�ti�?Pj S�l����WS�u�uj�u�օ�t�uPS�u��`�E�S�x����E�Y�u3�9]u��@�E9]u��@�E�u��3  Y���u3��G;EtSS�MQ�uP�u��3  ����;�t܉u�u�u�u�u�u��`��;�tV�vl��Y�Ǎe�_^[�M�3��b���Ë�U����u�M���n���u$�M��u �u�u�u�u�u�������}� t�M��ap��Ë�U��V�u����  �v�l���v��k���v��k���v��k���v��k���v��k���6��k���v ��k���v$��k���v(�k���v,�k���v0�k���v4�k���v�k���v8�k���v<�k����@�v@�k���vD�|k���vH�tk���vL�lk���vP�dk���vT�\k���vX�Tk���v\�Lk���v`�Dk���vd�<k���vh�4k���vl�,k���vp�$k���vt�k���vx�k���v|�k����@���   ��j�����   ��j�����   ��j�����   ��j�����   ��j�����   ��j�����   �j�����   �j�����   �j�����   �j�����   �j����,^]Ë�U��V�u��t5�;�tP�mj��Y�F;�tP�[j��Y�v;5�tV�Ij��Y^]Ë�U��V�u��t~�F;��tP�'j��Y�F;��tP�j��Y�F;��tP�j��Y�F; �tP��i��Y�F;�tP��i��Y�F ;�tP��i��Y�v$;5�tV�i��Y^]��������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U���S�u�M��k���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�/����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M���j���E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���58�N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�4���+8�;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�58�N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��<�A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;0��<���   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�0��D��3�@�   �D��e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+<���M���Ɂ�   �ً@�]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5P�N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�L���+P�;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5P�N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��T�A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;H��T���   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�H��\��3�@�   �\��e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+T���M���Ɂ�   �ًX�]���@u�M�U�Y��
�� u�M�_[�Ë�U���|���3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u����SSSSS�    聻����3��N  �U�U��< t<	t<
t<uB��0�B���/  �$��-�Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�a#  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �"  =�����.  �����`�E�;���  }�ع ��E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��K
3��E��EԉE؉E܋E΋��  3�#�#ʁ� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uB�E����u9u�u9u�u3�f�E���  f;�u!B�C���u9su93u�ủuȉu���  �u��}��E�   �E��M���M���~R�DĉE��C�E��E��M��	� �e� ���O��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?�����  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋M��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9M�w�Mԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�B�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�U�f�EċE؉EƋE܉E�f�U��3�f�����e� H%   � ���e� �Ẽ}� �<����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[�M���Ð�'�'/(b(�(�(�(N)9)�)�)\)��U���t���3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�f��t�C-��C �u�}�f��u/��u+��u'3�f;�����$ f��C�C�C0�S3�@�  ��  f;���   3�@f��   �;�u��t��   @uh���Qf��t��   �u��u;h���;�u0��u,h���CjP������3���tVVVVV蔲�����C�*h���CjP������3���tVVVVV�h������C3��q  �ʋ�i�M  �������Ck�M��������3���f�M๠��ۃ�`�E�f�U�u�}�M�����  }� ��ۃ�`�E�����  �E�T�˃������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE��P
3ɉM��M��M�M��M��3�� �  �u���  #�#֍4
����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��{����M�����?  ��  f;���  �E�3҉U��U��U�U��U��ɋ�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��V���3�3�f9u���H%   � ���E��\���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �^�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[��C���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95(���  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��{���Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��U��SVWUj j h\;�u�b!  ]_^[��]ËL$�A   �   t2�D$�H�3��@?��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�hd;d�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �yd;u�Q�R9Qu�   �SQ�`��SQ�`��L$�K�C�kUQPXY]Y[� ��������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ��U��j
j �u�  ��]�������Q�L$+ȃ����Y�*  Q�L$+ȃ����Y�  ��U��QQ�EV�u�E��EWV�E��  ���Y;�u蒕��� 	   �ǋ��J�u�M�Q�u�P��`�E�;�u�`��t	P脕��Y�ϋ�����@������D0� ��E��U�_^��jh���si������u܉u��E���u�)����  ����� 	   �Ƌ���   3�;�|;4�r!������8����� 	   WWWWW�H������ȋ�����@���������L1��u&辔���8褔��� 	   WWWWW������������[P�  Y�}���D0t�u�u�u�u�������E܉U���V���� 	   �^����8�M���M���E������   �E܋U��h����u�@  YË�U���  �g  ���3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�����0�ғ��VVVVV�    �5���������  SW�}�����4�@������ǊX$�����(�����'�����t��u0�M����u&胓��3��0�g���VVVVV�    �ʢ�����C  �@ tjj j �u�~������u�i  Y����  ��D���  �V���@l3�9H�������P��4�� �����`���`  3�9� ���t���P  ��`��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P�Z���Y��t:��4���+�M3�@;���  j��@���SP�[  �������  C��D����jS��@���P�7  �������  3�PPj�M�Qj��@���QP�����C��D�����`�����\  j ��<���PV�E�P��(���� �4��`���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4��`����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@����D  Yf;�@����h  ��8����� ��� t)jXP��@����  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4��`���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4��`���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  ��`��;���   j ��,���P��+�P��5����P��(���� �4��`��t�,���;����`��@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0��`��t��,�����@��� ��8�����`��@�����8��� ul��@��� t-j^9�@���u�Z���� 	   �b����0�?��@����f���Y�1��(�����D@t��4����8u3��$�����    �"����  ������8���+�0���_[�M�3�^�Y4����jh���'a���E���u�����  �ˌ��� 	   ����   3�;�|;4�r!轌���8裌��� 	   WWWWW�������ɋ�����@���������L1��t�P��  Y�}���D0t�u�u�u�.������E���@���� 	   �H����8�M���E������	   �E��`����u�1  YË�U��� �h   ��R��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u赋��� 	   3�]�V3�;�|;4�r藋��VVVVV� 	   �������3���ȃ�����@����D��@^]øp�á �Vj^��u�   �;�}�ƣ �jP�RR��YY�����ujV�5 ��9R��YY�����ujX^�3ҹp�������� �����|�j�^3ҹ��W������@�����������t;�t��u�1�� B���|�_3�^��  �=�� t��  �5���;��YË�U��V�u�p�;�r"��вw��+�����Q�)���N �  Y�
�� V��`^]Ë�U��E��}��P��~���E�H �  Y]ËE�� P��`]Ë�U��E�p�;�r=вw�`���+�����P��}��Y]Ã� P��`]Ë�U��M���E}�`�����Q�}��Y]Ã� P��`]Ë�U��EV3�;�u蚉��VVVVV�    ������������@^]á����3�9$�����Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�$���j^SSSSS�0舘�������V�u�M��<���E�9X��   f�E��   f;�v6;�t;�vWSV�9�����ш��� *   �ƈ��� 8]�t�M��ap�_^[��;�t2;�w,覈��j"^SSSSS�0�
�����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p��`;�t9]�^����M;�t����`��z�D���;��g���;��_���WSV�8�����O�����U��j �u�u�u�u�|�����]Ë�U������3ŉE�j�E�Ph  �u�E� ��`��u����
�E�P����Y�M�3��/���Ë�U���4���3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5�`�M�QP�֋�`��t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��4�����YF;�~[�����wS�D6=   w/������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�6��Y;�t	� ��  ���E���}�9}�t؍6PW�u��<7����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u��`��t`�]��[��`9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�NM��YY�E�;�t+WWVPV�u�W�u��;�u�u��07��Y�}���}��t�MЉ�u�衬��Y�E��e�_^[�M�3��M-���Ë�U������3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[�+���Ë�U���VW�u�M��7���E�u3�;�t�0;�u,����WWWWW�    �I������}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�����M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&�E����E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9x�uhЭ�P������]����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ���U��MS3�;�VW|[;4�sS������<�@��������@t5�8�t0�=L�u+�tItIuSj��Sj��Sj�� a���3������� 	   ��������_^[]Ë�U��E���u������  �ހ��� 	   ���]�V3�;�|";4�s�ȃ�����@�����@u$踀���0螀��VVVVV� 	   ����������� ^]�jh���T���}����������4�@��E�   3�9^u6j
�u��Y�]�9^uh�  �FP����YY��u�]��F�E������0   9]�t����������@��D8P��`�E��|T���3ۋ}j
��s��YË�U��E�ȃ�����@����DP��`]Ë�U������3ŉE�V3�95`�tO�=Զ�u�g  �Զ���u���  �pV�M�Qj�MQP�a��ug�=`�u��`��xuω5`�VVj�E�Pj�EPV�aP��`�Զ���t�V�U�RP�E�PQ�a��t�f�E�M�3�^�n&�����`�   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��m2���E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�G���YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p��`���E�u�M;��   r 8^t���   8]��e����M��ap��Y����~��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p��`���:���뺋�U��j �u�u�u�������]�jh����Q��3ۉ]�j�sr��Y�]�j_�}�;= �}W��������9tD� �@�tP�  Y���t�E��|(������ P�l`����4�p.��Y����G��E������	   �E��Q���j�q��YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�C���YP�������;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�����P�  Y��Y��3�^]�jh ��P��3��}�}�j�!q��Y�}�3��u�;5 ���   �����98t^� �@�tVPV�����YY3�B�U�������H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u����4�V�����YY��E������   �}�E�t�E��1P���j�o��Y�j����Y����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h��a�ԶáԶV�5a���t���tP�֡ж���t���tP��^Ë�U��SV�uW3����;�u��z��WWWWW�    �&�������B�F�t7V�{���V����  V�����P�   ����}�����F;�t
P�+��Y�~�~��_^[]�jh(��N���M��3��u3�;���;�u�@z���    WWWWW裉���������F@t�~�E��N���V����Y�}�V�*���Y�E��E������   �ՋuV�����Y�jhH��$N���E���u��y��� 	   ����   3�;�|;4�r�y��� 	   SSSSS�������Ћ����<�@���������L��t�P�����Y�]���Dt1�u�g���YP�a��u�`�E���]�9]�t�Ny���M��1y��� 	   �M���E������	   �E��M����u�)���YË�U��V�uWV� ���Y���tP�@���u	���   u��u�@Dtj�����j�������YY;�tV�����YP�a��u
�`���3�V����������@�����Y�D0 ��tW�x��Y����3�_^]�jhh��L���E���u�fx���  �Kx��� 	   ����   3�;�|;4�r!�=x���8�#x��� 	   WWWWW膇�����ɋ�����@���������L1��t�P�g���Y�}���D0t�u�����Y�E����w��� 	   �M���E������	   �E��6L����u�����YË�U��V�u�F��t�t�v�(���f����3�Y��F�F^]�����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%�`������������h�\�U)��Y����̃=� uK� ���t���Q<P�B�Ѓ�� �    ����tV���`F��V躎������    ^�                                                                                                                                                                                                           ̋ �  � � � .� :� L� `� t� �� ��  ֌ � �� � � � 4� D� \� d� r� �� �� �� �� ̍ � �� � .� D� ^� l� z� �� �� �� Ȏ � � � � .� <� H� T� ^� j� |� �� �� �� ҏ � � 
� � ,� >� P� `� r� �� �� �� �� Ɛ Ԑ         �\        Ԫ��R��G        PX�H                <0N       p   �� �u bad allocation                    �?    USERNAME         @�@ikto    ikfrom  texturesearchpath   dst src fbx c4d c:\buildagent\work\b2b44f52c74c2f2a\src\source\convert.cpp  EXPORT_ERROR: An unknown error has occured  EXPORT_ERROR: An error occured while saving the document    EXPORT_ERROR: Destination bad format    EXPORT_ERROR: Source bad format EXPORT_ERROR: Source either does not exist or cannot be located EXPORT_ERROR: An error occured while loading the document   EXPORT_ERROR: FBX exporter not found    SUCCESS framerate=  version=    -UnityC4DFBXtmp -UnityC4DFBXout 0   Filtered:       Name: ' '   Plugin:     Processing  Scanning    -UnityC4DFBXcmd * (c) 2006-2011 Unity Technologies ApS - http://unity3d.com * Unity-C4DToFBXConverter for Cinema 4D R12. Version: 3.09  ����MbP?D��� �k ��`�     c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_baseobject.cpp c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_general.h  %s     c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_file.cpp       c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_basetime.cpp             �? �Ngm��C   ����A  4&�k�  4&�kC؄p� c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_resource.cpp   #   M_EDITOR        �������������c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_libs\lib_ngon.cpp  c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_pmain.cpp  res     c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_basebitmap.cpp  ��y    c:\buildagent\work\b2b44f52c74c2f2a\sdk\r12\_api\c4d_gv\ge_mtools.cpp   h��y��py�� z�z��    D��}      �?      �?3      3            �      0C       �       ��              e+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    P���EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:                �������             ��      �@      �              �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow       �?5�h!���>@�������             ��      �@      �            	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        hv`vTvHv<v0v$vvvv�aHq,qq�p�p�u�u�p�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u�u|uxutupuluhudu`u\uXuTuHu<u4u(uuu�t�t�t�tptPt,tt�s�s�s�sxstsls\s8s0s$ss�r�r�r�r`r4rr�q�q�qxq\q�aGetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun 1#QNAN  1#INF   1#IND   1#SNAN  SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           ����   RSDSBbQۻt�C�UO��NT�   C:\BuildAgent\work\b2b44f52c74c2f2a\src\obj\Unity-C4DToFBXConverter12_Win32_Release.pdb             �(�    l�        ����    @   �            ��X�           h�p�    ��        ����    @   X�            ����           ����(�    ��       ����    @   ��            ܠ�           ���    ܠ        ����    @   �            ,�4�           D�L�    ,�        ����    @   4�            H�|�           ����    H�        ����    @   |�            h�ą           ԅ��(�    h�       ����    @   ą            ���            �(�    ��        ����    @   �            ġX�           h�p�    ġ        ����    @   X�     � d� d;                     ����    ����    �����|�|    ����    ����    ����    '�    ����    ����    ����    Є    ����    ����    ����    )�    ����    ����    ����    [�����    j�����    ����    ����    �����    )�����    ����    ����    ��    ����    ����    ����_�c�    ����    ����    ����?�[�    ����    ����    ����    H�    ����    ����    ����    �    ����    ����    ����    Q�    ����    ����    ����    K�    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    X�    ����    ����    ����[�o�    ����    ����    ��������    ����    ����    ����    ��    ����    ����    ����(�?�    ����    ����    ����0L    ����    ����    ����    0?    ����    ����    ����    ?G    ����    ����    ����    jS    ����    ����    ����    +V    ����    ����    ����    �W        �W����    ����    ����    eY    ����    ����    ����    GZ    ����    ����    ����    �[��         ܋  `                     ̋ �  � � � .� :� L� `� t� �� ��  ֌ � �� � � � 4� D� \� d� r� �� �� �� �� ̍ � �� � .� D� ^� l� z� �� �� �� Ȏ � � � � .� <� H� T� ^� j� |� �� �� �� ҏ � � 
� � ,� >� P� `� r� �� �� �� �� Ɛ Ԑ     ZGetTempPathA  KERNEL32.dll  �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �GetLastError  �HeapFree   GetProcAddress  �GetModuleHandleA  -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent �GetModuleHandleW  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �InterlockedIncrement  �SetLastError  �InterlockedDecrement  !Sleep ExitProcess �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA � DeleteCriticalSection �GetModuleFileNameA  JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW zWideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy WVirtualFree TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �WriteFile �LeaveCriticalSection  � EnterCriticalSection  TVirtualAlloc  �HeapReAlloc �HeapSize  [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �LoadLibraryA  �InitializeCriticalSectionAndSpinCount �RtlUnwind �GetLocaleInfoA  ZRaiseException  �LCMapStringA  MultiByteToWideChar �LCMapStringW  =GetStringTypeA  @GetStringTypeW  �SetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW x CreateFileA C CloseHandle AFlushFileBuffers              <0N    "�          � �  � p, @�   Unity-C4DToFBXConverter12.cdl c4d_main                                                                                                                                                                                        |a    |a    B�     b�     a�     `�     ��    ��    qr            |a|a|a|a|a|a|a�g    .?AVGeSortAndSearch@@   �g    .?AVNeighbor@@  �g    .?AVDisjointNgonMesh@@  |a|a|a|a|a|a�g    .?AVBaseData@@  |a|a|a|a|a|a|a|a|a|a|a|a|a|a�g    .?AVGeToolNode2D@@  �g    .?AVGeToolDynArray@@    �g    .?AVGeToolDynArraySort@@    �g    .?AVGeToolList2D@@  |au�  s�  N�@���D    |a�g    .?AVtype_info@@     fmod         ��V��V���V��V�����V�V��V�sqrt    ��������������������    �����
                                                                   x   
   |a                  �n   Tn	   (n
   �m   dm   4m   m   �l   �l   �l   Ll   l   �k   �k   hk    0k!   8j"   �ix   �iy   tiz   di�   `i�   Pi       ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ���������������ƶ̶Ҷ��	��*�:�N�^�~�������·ַ��"�'�A�F�f�z�����Ƹ˸��
��6�J�j�o�������¹ڹ���-�2�R�f�~�������Ѻֺ��
�"�  ?                                                                                                                                                                                                                                                                                                                         	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                                                                             abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     ���  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    \|����C                                                                                              �            �            �            �            �                              �        Xz�~`�(��   ���        xxhx�&         p   p   �o    p   Ly   Dy!   <y   �o   �o   �o   4y   ,y   �o   �o    �o   �o   �o   $y   �o   y   y   y   y   �x"   �x#   �x$   �x%   �x&   �x      �      ���������              �       �D        � 0     XzZ|    ������|�x�t�p�h�`�X�L�@�8�,�(�$� �������� �������؁�Ёȁ����������������l�`�	         (�.   �����������   .                 ���5      @   �  �   ����              �             �     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �p     ����    PST                                                             PDT                                                              �@�����        ����                 �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
       ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l      ��������                                                                                                                                                                                                                                                                                                             0"000A0N0d0�0�0�0�01'151D1t1�1�1�1�1�122�2�2�2b3�3�3�3444K4]4o4�4�4�4�4�4�4�45:5\5�5�56:6v6�6�6�67-7K7i7�7�7;8W8p8�8�89�9�9�9�9�9
:,:>:P:�:�:�:�:�:�:;!;3;?;N;g;�;�;�;�;�;�;
<<-<M<[<q<�<�<�<�<�<==*=J=d=x=�=�=�=�=�=>>e>�>�>�>�>�>9?�?�?�?      4  	040P0j0�0�0�0�001�1�12)2]2�2�2�2�2,3>3O3a3s3�3�3�3�3�3(4:4L4]4�4W5l5�5�5�5�5�5�5�56&6;6O6a6v6�6�6�6�6�6�67:7Z7x7�7�7�7�78$858G8P8e8z8�8�8�8�8�8�8�829�9�9�9�9�9�9 ::A:R:d:m::�:�:�:�:�:�:�:�:;;';=;O;X;i;{;�;<<0<L<a<|<�<�<�<=%=:=B=[=z=�=�=�=�=�=>6>;>P>e>n>�>�>�>�>�>??,?5?K?�?�?�?�?�?�?   0  <  00!060J0\0n0w0�0�0�0�0�0111P1e1v1�1�1�1�1�12222222 2$2(2,202a2s2�2�2�2�2�2�2�2�2313G3[3r3�3�3�3�3�3�34&4B4X4k4~4�4�4�4�4�455&585J5[5�5�5�5�5�5�566)626D6V6~6�6�6�6�6�6�6737E7V7h7�7�7�7�7�7�78]8|8�8�8�8 99#959G9r9�9�9�9�9�9�9$:D:d:v:�:�:�:�:; ;2;C;U;g;x;�;�;<<�<=B=u=�=�=%>u>�>�>?E?�?�? @  �   0_0�0�0"1R1�1�12b2�2�2"3U3�3�3454e4�45E5�5�56#6P6d6t6�6�6%7e7�7�758u8�8999a9�9�9�9�9�9:::e:�:�:�:(;O;�;�;�;5<]<�<�<�<"=V=x=�=U>r>�>�>�>�>?$?D?a?q?�?�?�?�?�?�?   P  �   040T0t0�0�0�0�01D1d1�1�1�1�12$2D2�2�2�2�2�23!3?3a33�3�3�3414T4t4�4�4�4�45$5A5T5t5�5�5�5646a6�6�6�67d7�7�7848T8t8�8�8�8�8$949d9�9�9�9:$:Q:t:�:�:�:!;D;�;�;�;�;<1<Q<q<�<�<�<�<=1=Q=q=�=�=�=�=>D>d>�>�>�>?$?A?d?�?�?�?   `  �   040d0�0�0�0B1a1�1�1�1�12A2a2�2�2�2�23D3t3�3�3�34$4D4q4�4�4�4�45 5D5�5616D6d6�6�6�6717a7�7�7�7�7848�8�8�8�8$9T9t9�9�9*:k:�:�:�:;$;T;�;�;�;�;�;�;:<T<�<�<�<=d=�=�=b>�>?%?:?]?�?�?�? p  �   060_0�0�0�01H1y1 2D2T2�2�2�2	333G3e3�3�3�3�34D4d4�4�4�4�45a5�5�5�56!6D6d6�6�6�6$7q7�7�7�7�7?8^8z8�8�8�8(9C9q9�9�9�9�9:&:V:x:�:�:�:�:;3;H;�;�;�;�;<+<K<`<|<7=J=�=�=�=�=>L>   �  �   [0
3#3t3�3�3�34D4_4666 6�6�6�6�6�6!747d7�7�7�7�7$8T8t8�8�89$9T9t9�9�9�9�9:4:F:a:t:�:�:�:�:�:;4;q;�;�;�;�;<4<T<q<�<�<�<�<�<=$=D=d=�=�=�=�=>1>D>d>�>�>�>�>?T?z?�?�?�?   �  �   0$0D0d0�0�0�0�01D1�1�1�1C2�2�2�23D3q3�3�3�3�34!444T4t4�4�4�4	55r5�5�5�56$6D6�6�6�6�6�67&767d7�7�7�7�7808D8T8t8�8�8�8
9=9K9^9s9�9�9�9�9�9:":2:T:x:�:�:�:�:%;S;i;w;�;�;�;�;#<9<G<V<�<�<�<�<$=M={=�=�=�=>/>T>t>�>�>�>�>?$?D?a?t?�?�?�?   �  (  040T0t0�0�0�0�01!141Q1d1�1�1�1�1�12%262H2d2�2�2�2�2�233#3D3U3c3�3�3�3�3�34!4D4\4p4�4�4�4�4�4�45 5D5\5p55�5�5�5�56!646T6t6�6�6�6�67747d7�7�7�7�78$8Q8d8�8�8�8�89$9D9a9q9�9�9�9�9�9:4:T:t:�:�:�:;;/;P;X;l;�;<;<Q<u<�<�<�<=4=T=t=�=�=�=�=>4>Q>a>t>�>�>�>�>�>�>?4?S?a?p?�?�?�?   �  ,  00!010A0Q0d0�0�0�0�0�0�01$1D1d1�1�1�1�12$2W2p2�2�2�2�2�23'393d3�3�3�3�34$4;4O4^4n4�4�4�4�4�4�45$5H5n5�5�5�5�5�5�56646R6f6u6�6�6�6�6$717A7T7t7�7�7�7�7848T8t8�8�8�8�8949T9t9�9�9�9�9:4:\:�:�:�:�:;4;T;t;�;�;�;�;<4<T<t<�<�<�<�<=4=T=t=�=�=�=�=>$>D>d>�>�>�>�>�>�>?$?D?f?z?�?�?�?�?   �  �   00-0`0u0�0�0141Q1d1�1�1�1�12D2t2�2�2�2�23$3Q3d3�3�3�3�3424Q4t4�4�4�4$5D5a5�5�5�5�56D6q6�6�6�67A7a7�7�7�7�78$8D8d8�8�8�8�8�8949T9�9�9�9l:�:�:;q;�;
<-<�<�<�<a=~=�=>.>C>�>�>?A?d?�?   �  �   S0|0�0#1L1t1�12D2�2�2�2k3�34a4�4�45a5�5�5L6�6�67�7�7�7>8^8s8�8!9�9�9$:D:a:q:�:�:�:�:;4;d;�;�;�;<$<D<a<�<�<�<=0=R=�=�=�=�=>&>a>�>�>�>�>?�?�?�?�?�?�? �  �   0D0a0t0�0�0�01D1d1�1�1�1�1�1'2b2�2�2�223`3�3�344G4g4�475u5�5�5�5�5686V6d6�6�6$727Q7a7t7�7�7�78848T8|8�8�8�8$9D9a9�9�9I:e:�:�:I;e;�;�;<,<H<d<�<�<=%=�=�=!>�>�>�>�>?$?1?_?�?�?�?�?   �  @  0*080G0{0�0�01;1v1�1�1�1�1�122262I2[2m22�2�2�2�2�23$353H3t3�3�3�3�3�3�3�3�3444F4b4x4�4�4�4�4�4 5525C5V5�5�5�5�5�5�5�5�56&6D6V6r6�6�6�6�6�6�67&7B7T7f7o7�7�7�7�78"8/8G8Y8k8}8�8�8�8�8�89949F9X9a99�9�9�9�9�9�9:>:T:r::�:�:�:�:�:';T;q;�;<
<<&<0<K<g<�<�<�<�<�<=F=h=�=�=>>!>4>�>�>�>�>�>
??B?_?�?�?   @   D0Y0{0�0�1�1�12$2D2d2�2�2�2�2343T3t3�3�3�3414�4�4??    D   !9A9m9�9�9%:u:�:�:2;b;�;�;<E<�<�<=B=r=�=�=>5>u>�>?U?�?�?   �   0U0�01e1H3i3�5h6l6p6t6x6[7i7�7�7"808U8]89,9P9^9�9�9�:�:�:�:`;n;�;�;R<X<�<�<�<�<�<�<�<2=E=_=x=|=�=�=�=�=�=�=�=%>k>�>5?u?�? 0 �   0F0�0�01H1�1�1%2e2�2353x3�34B4u4�4�45e5�5�5�56*6R6�6�6%7r7�78U8�8�8E9�9�9:R:�:�:(;�;�;(<�<�<%=v=�=>e>�>?H?�?   @ t   H0�01E1�1�12e2�2�2E3�3�324u4�45f5�56U6�6�6�67e7�7�758�8�8%9�9�96:�:�:;E;�;�;<e<�<=5=�=�=>4>|>�>/?�? P �   ,0t0�0�0�0�0!1d1�1�1f2�2]3�3#4Q4n4�4�446�6�6�7�78D8�8�8�8949T9�9�9�9M:x:�:�:�:�:�:�:�:�:;;; ;';.;5;<;C;J;Q;X;_;j;�;�;�;�<%=�>�>?$?A?T?�?�?�?�? ` �   040T0�0�0�0�0$1D1d1�1�122'2d2�2�2�23!3D3d3�3�3�3�3!4�4�4�4$5A5T5(7:7M7p7(9a9t9�9�9�9!:1:S:t:�:�:�:;7;E;T;�;�;�;�;�;$<T<8=l=�=�=;>??&?�?�?�?   p �   B0�0�0141e1�12W2h2:6�6�68@8�8�8�8�89&9M9�9�9B:G:M:Q:W:[:a:e:k:o:t:z:~:�:�:�:�:�:�:�:�:;;;N;f;n;t;�;�;�;<'<?<�<�<2=N=�=:>o>�>�>�>�>�>�>�>�>??? ?$?(?,?0?4?~?�?�?�?�?�? � �   00#0(0,000Q0{0�0�0�0�0�0�0�0�0�01 1$1(1,1�1�1�1�1
2#2�2�2�2�2�2�2F3L3l3�3�3 4}4�4�4�4�455�5�5�5�5�5�6�6�6�6�647<7Q7\7:�:�: � �  0�0t2�2�2�2�233+31373=3C3I3P3W3^3e3l3s3z3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3444-434>4J4_4f4z4�4�4�4�4�4�4�4�4�45 5&525A5G5P5\5j5p5|5�5�5�5�5�5�5�5�5�5696y66�6�6�6�6	7�7�7�7�7�7<8L8R8^8d8t8z8�8�8�8�8�8�8�8�8�8�8�8�8�89999(9-92989<9B9G9M9R9a9w9�9�9�9�9�9�9�9�9�9�9�9�9:J:S:_:�:�:�:�:�:�:;&;S;n;t;};�;�;<< <+<0<@<J<Q<\<e<{<�<�<�<�<�<�<=&=P=U=`=e=�=>>%>9>Z>`>�>�>�>1?;?c?|?�?�?�?   � �   Q0W0{0�0�0�0�011g1r1|1�1�1K3\3d3j3o3u3�3�3�344+484?4v4�4�4
5#52575X5]5�5�5�5�5�5�5�5�5�5�5�56666:6�6�6�6�6�7�78�8�89$9{9�9�9�9�9�9�9�9::%:�:�:;	;�;�;"<�<�<=M=e=p=�=�=�=�=�=�=>?>d>w>�>�>�>�> � <   D1�1�1�2�2�2�2�2�2�3@4�4\5�5�5�566x6�6�=�>?U?�?   � �    0"0]0�1�12�2�2�2;3C3P3�3�34&4A4M4Y4e4�4�4�4�4�4�4�4�45555*565?5H5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5B6�6�6�6�6�6�67$7=7Q7W7`7s7�7,8L8Z8_8�:�:�:�:�:�:�:�:;;*;5;;;A;F;O;l;r;};�;�;�;�;�;�;�;�;�;�;�;�;�;�;<#<)<:<�<   � �   ;0G0z0�0�01�2�23$3@3c3v3�3�3�4�4=5C5677-757E7V7�7,8C8�9�9:::&:/:9:m:x:�:�:�:�:�:;H;[;�;�;0<�<�<0=<=O=a=|=�=�=�=�=�=�=�=�=�=>+>T>e>�>M?w?�? � �   0]0�01"131o1�1�1�2�2�2�2�2�2J3V3�4�4c5:6o6�6�6�6�6�6�6�6�6777 7$7(7,70747~7�7�7�7�7�788#8(8,808Q8{8�8�8�8�8�8�8�8�8�89 9$9(9,9�;�=�=[>p>�>�>�>?P?�?�?�? � �   J0P0t0�0�0�0�0$1�1�1�12!2'2�2�2�2�2�2�2�2�2.3<3�3�3�3�3�3�3�3�3Y4b4h4�45
55O5�5�57=7K7Q7a7f7~7�7�7�7�7�7�7�7�7�7�7�718N8k8�9�9�9(;/;:<�<�< =�=�=�=     @   �0�1s3�3�3�5�7�7�7�7�7�7�7�7�7�8.;�<�<�<�<�<N=W>�>�>]?�?  h   �1�1�122!2Q2~2�2�2�2�2�2�2�2&3�3m4�45�5g6q6�6�6�6�6�6�6�67�7::%:G:Y:k:}:�:�:�:�<�=�=�>r?     \   00�0�0�0i1�1#23!3�3�4O5U5�5�56�6�6�6�7Q:h:�=�=�=�=�=�=�=�=�=�=�=�=�=�>�>�>?z?�? 0 (   �9P;�;�;9<S<\<�=�=>$>b>�>J?�?   @ p   c0�0s1�1�1�3c4,5]5s5�5�5p6�6�6P7�7�7�7�78&838?8O8V8e8q8~8�8�8�8�8�89:9I9R9v9�9�9�9;2;�;�;�;<<�<=�= P �   �1�1�1�1292�2�2�2�2R3]3�3�3�3�3�3�3�3�3�344#4)4?4Z4�4m5�5�5�5�5�5�56�6
7787�7@8F8K8Q8X8j8�8s9�9�9�9:h:�:�:�:�:$;S;�<�<�<�<�<==+= ` D   $1014181<1@1L1P1�4�4�4�4�4�5�5,707�7�7�7�7�7�7�7�7�7�7�7@8D8 p �   x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 � �   �3�34 4(4@4P4T4d4h4p4�4�4�4�4�4�4�4�4�4�4�4�455,505@5D5L5d5t5x5�5�5�5�5�5�5�5�5�5�5�5666 6(6@6P6T6d6h6p6�6�6�6�67(7H7T7p7|7�7�7�7�7�7�7888X8x8�8�8�8�8�89989T9X9t9x9�9�9�9�9:$:@:`:�: �    00P0T0X0\0`0d0h0l0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1H1h1�1�1�1�1�1�1�1�1 22222222 2$2(2,282<2@2D2H2L2P2T2X2\2h2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�34"4&4*4.42464:4>4B4F4J4N4R4V4Z4^4b4f4j4n4r4v4z4~4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�455
55555�;�<H=X=h=x=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>? ?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   �     00000p0x0�3�3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  